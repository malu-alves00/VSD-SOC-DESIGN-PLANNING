module picorv32a (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 sky130_fd_sc_hd__nand2_1 _21192_ (.A(net237),
    .B(net521),
    .Y(_18523_));
 sky130_fd_sc_hd__nor2_4 _21193_ (.A(mem_do_wdata),
    .B(mem_do_rdata),
    .Y(_18524_));
 sky130_vsdinv _21194_ (.A(mem_do_rinst),
    .Y(_18525_));
 sky130_fd_sc_hd__o21ai_2 _21195_ (.A1(_18523_),
    .A2(_18524_),
    .B1(_18525_),
    .Y(_18526_));
 sky130_fd_sc_hd__buf_2 _21196_ (.A(_18523_),
    .X(_18527_));
 sky130_fd_sc_hd__nand2_1 _21197_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_18528_));
 sky130_fd_sc_hd__nor2_8 _21198_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_00290_));
 sky130_fd_sc_hd__a21oi_2 _21199_ (.A1(_18527_),
    .A2(_18528_),
    .B1(_00290_),
    .Y(_18529_));
 sky130_fd_sc_hd__nand2_4 _21200_ (.A(_18526_),
    .B(_18529_),
    .Y(_18530_));
 sky130_vsdinv _21201_ (.A(net101),
    .Y(_18531_));
 sky130_fd_sc_hd__buf_6 _21202_ (.A(_18531_),
    .X(_18532_));
 sky130_fd_sc_hd__clkbuf_4 _21203_ (.A(_18532_),
    .X(_18533_));
 sky130_fd_sc_hd__a21oi_2 _21204_ (.A1(_18530_),
    .A2(mem_do_prefetch),
    .B1(_18533_),
    .Y(_18534_));
 sky130_vsdinv _21205_ (.A(mem_do_rdata),
    .Y(_18535_));
 sky130_vsdinv _21206_ (.A(\cpu_state[6] ),
    .Y(_18536_));
 sky130_fd_sc_hd__nor2_1 _21207_ (.A(_18535_),
    .B(_18536_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _21208_ (.A(_18534_),
    .B(_00319_),
    .Y(_18537_));
 sky130_vsdinv _21209_ (.A(_18537_),
    .Y(_18538_));
 sky130_fd_sc_hd__nor2_2 _21210_ (.A(_00332_),
    .B(_18538_),
    .Y(_18539_));
 sky130_fd_sc_hd__clkbuf_2 _21211_ (.A(net101),
    .X(_18540_));
 sky130_fd_sc_hd__buf_2 _21212_ (.A(_18540_),
    .X(_18541_));
 sky130_fd_sc_hd__clkbuf_4 _21213_ (.A(_18541_),
    .X(_18542_));
 sky130_fd_sc_hd__clkbuf_4 _21214_ (.A(_18542_),
    .X(_18543_));
 sky130_fd_sc_hd__buf_2 _21215_ (.A(\cpu_state[6] ),
    .X(_18544_));
 sky130_vsdinv _21216_ (.A(_18539_),
    .Y(_18545_));
 sky130_fd_sc_hd__a21o_1 _21217_ (.A1(instr_lb),
    .A2(_18544_),
    .B1(_18545_),
    .X(_18546_));
 sky130_fd_sc_hd__o211a_1 _21218_ (.A1(latched_is_lb),
    .A2(_18539_),
    .B1(_18543_),
    .C1(_18546_),
    .X(_04071_));
 sky130_fd_sc_hd__buf_2 _21219_ (.A(_18540_),
    .X(_18547_));
 sky130_fd_sc_hd__buf_2 _21220_ (.A(_18547_),
    .X(_18548_));
 sky130_fd_sc_hd__clkbuf_4 _21221_ (.A(_18548_),
    .X(_18549_));
 sky130_fd_sc_hd__a21o_1 _21222_ (.A1(instr_lh),
    .A2(_18544_),
    .B1(_18545_),
    .X(_18550_));
 sky130_fd_sc_hd__o211a_1 _21223_ (.A1(latched_is_lh),
    .A2(_18539_),
    .B1(_18549_),
    .C1(_18550_),
    .X(_04070_));
 sky130_vsdinv _21224_ (.A(instr_retirq),
    .Y(_18551_));
 sky130_fd_sc_hd__nand2_1 _21225_ (.A(_18551_),
    .B(net518),
    .Y(_18552_));
 sky130_vsdinv _21226_ (.A(_00331_),
    .Y(_18553_));
 sky130_fd_sc_hd__nand2_1 _21227_ (.A(_18552_),
    .B(_18553_),
    .Y(_18554_));
 sky130_vsdinv _21228_ (.A(latched_branch),
    .Y(_18555_));
 sky130_fd_sc_hd__nand2_1 _21229_ (.A(_18554_),
    .B(_18555_),
    .Y(_18556_));
 sky130_fd_sc_hd__o211a_1 _21230_ (.A1(_21141_),
    .A2(_18554_),
    .B1(_18549_),
    .C1(_18556_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_4 _21231_ (.A(_18533_),
    .X(_18557_));
 sky130_fd_sc_hd__nand2_1 _21232_ (.A(\mem_state[0] ),
    .B(mem_do_rinst),
    .Y(_18558_));
 sky130_fd_sc_hd__o211a_1 _21233_ (.A1(\mem_state[0] ),
    .A2(_18527_),
    .B1(\mem_state[1] ),
    .C1(_18558_),
    .X(_18559_));
 sky130_vsdinv _21234_ (.A(_00290_),
    .Y(_18560_));
 sky130_fd_sc_hd__nor2_1 _21235_ (.A(mem_do_rinst),
    .B(mem_do_prefetch),
    .Y(_18561_));
 sky130_vsdinv _21236_ (.A(_18561_),
    .Y(_18562_));
 sky130_fd_sc_hd__nor2_1 _21237_ (.A(mem_do_rdata),
    .B(_18562_),
    .Y(_18563_));
 sky130_fd_sc_hd__inv_2 _21238_ (.A(mem_do_wdata),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_2 _21239_ (.A(_18563_),
    .B(_00291_),
    .Y(_18564_));
 sky130_fd_sc_hd__nor2_1 _21240_ (.A(_18560_),
    .B(_18564_),
    .Y(_18565_));
 sky130_fd_sc_hd__nor3_2 _21241_ (.A(net408),
    .B(_18559_),
    .C(_18565_),
    .Y(_18566_));
 sky130_fd_sc_hd__o21a_1 _21242_ (.A1(_18557_),
    .A2(_18566_),
    .B1(_00300_),
    .X(_18567_));
 sky130_fd_sc_hd__nor2_2 _21243_ (.A(net408),
    .B(_18557_),
    .Y(_18568_));
 sky130_fd_sc_hd__clkbuf_2 _21244_ (.A(_18568_),
    .X(_18569_));
 sky130_fd_sc_hd__and2b_1 _21245_ (.A_N(_18567_),
    .B(\mem_state[1] ),
    .X(_18570_));
 sky130_fd_sc_hd__a31o_1 _21246_ (.A1(_21106_),
    .A2(_18567_),
    .A3(_18569_),
    .B1(_18570_),
    .X(_04068_));
 sky130_vsdinv _21247_ (.A(\mem_state[0] ),
    .Y(_18571_));
 sky130_fd_sc_hd__nor2_1 _21248_ (.A(_18571_),
    .B(_18567_),
    .Y(_18572_));
 sky130_fd_sc_hd__a31o_1 _21249_ (.A1(_21105_),
    .A2(_18567_),
    .A3(_18569_),
    .B1(_18572_),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_8 _21250_ (.A(_18532_),
    .B(_18530_),
    .Y(_18573_));
 sky130_vsdinv _21251_ (.A(_18573_),
    .Y(_18574_));
 sky130_fd_sc_hd__nor2_2 _21252_ (.A(_18525_),
    .B(_18574_),
    .Y(_18575_));
 sky130_fd_sc_hd__clkbuf_2 _21253_ (.A(_18575_),
    .X(_18576_));
 sky130_fd_sc_hd__buf_2 _21254_ (.A(_18576_),
    .X(_21108_));
 sky130_fd_sc_hd__inv_2 _21255_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_fd_sc_hd__clkbuf_2 _21256_ (.A(_18575_),
    .X(_18577_));
 sky130_fd_sc_hd__clkbuf_2 _21257_ (.A(_18577_),
    .X(_18578_));
 sky130_vsdinv _21258_ (.A(_00327_),
    .Y(_18579_));
 sky130_fd_sc_hd__or3_2 _21259_ (.A(\mem_rdata_latched[28] ),
    .B(_00330_),
    .C(_18579_),
    .X(_18580_));
 sky130_fd_sc_hd__and3b_1 _21260_ (.A_N(_00326_),
    .B(_00325_),
    .C(_00324_),
    .X(_18581_));
 sky130_fd_sc_hd__or4b_4 _21261_ (.A(_00329_),
    .B(_00328_),
    .C(_18580_),
    .D_N(_18581_),
    .X(_18582_));
 sky130_fd_sc_hd__nor2_1 _21262_ (.A(\mem_rdata_latched[27] ),
    .B(_18582_),
    .Y(_18583_));
 sky130_vsdinv _21263_ (.A(\mem_rdata_latched[25] ),
    .Y(_18584_));
 sky130_fd_sc_hd__nor3_2 _21264_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .Y(_18585_));
 sky130_fd_sc_hd__and4_1 _21265_ (.A(_18583_),
    .B(\mem_rdata_latched[26] ),
    .C(_18584_),
    .D(_18585_),
    .X(_18586_));
 sky130_fd_sc_hd__clkbuf_2 _21266_ (.A(_18586_),
    .X(_18587_));
 sky130_fd_sc_hd__nand2_1 _21267_ (.A(_18587_),
    .B(_18576_),
    .Y(_18588_));
 sky130_fd_sc_hd__or3b_1 _21268_ (.A(\mem_rdata_latched[26] ),
    .B(\mem_rdata_latched[25] ),
    .C_N(_18585_),
    .X(_18589_));
 sky130_fd_sc_hd__and2b_1 _21269_ (.A_N(_18589_),
    .B(_18583_),
    .X(_18590_));
 sky130_fd_sc_hd__o21ai_1 _21270_ (.A1(\mem_rdata_latched[19] ),
    .A2(_18590_),
    .B1(_18578_),
    .Y(_18591_));
 sky130_fd_sc_hd__o211ai_1 _21271_ (.A1(_00366_),
    .A2(_18578_),
    .B1(_18588_),
    .C1(_18591_),
    .Y(_04066_));
 sky130_fd_sc_hd__buf_2 _21272_ (.A(decoder_trigger),
    .X(_18592_));
 sky130_fd_sc_hd__nand2_1 _21273_ (.A(\cpu_state[1] ),
    .B(_18592_),
    .Y(_18593_));
 sky130_vsdinv _21274_ (.A(decoder_trigger),
    .Y(_18594_));
 sky130_vsdinv _21275_ (.A(\irq_mask[2] ),
    .Y(_18595_));
 sky130_vsdinv _21276_ (.A(\irq_pending[0] ),
    .Y(_18596_));
 sky130_fd_sc_hd__nor2_4 _21277_ (.A(\irq_mask[0] ),
    .B(_18596_),
    .Y(_18597_));
 sky130_vsdinv _21278_ (.A(\irq_pending[1] ),
    .Y(_18598_));
 sky130_fd_sc_hd__nor2_4 _21279_ (.A(\irq_mask[1] ),
    .B(_18598_),
    .Y(_18599_));
 sky130_vsdinv _21280_ (.A(\irq_mask[3] ),
    .Y(_18600_));
 sky130_fd_sc_hd__and2_1 _21281_ (.A(_18600_),
    .B(\irq_pending[3] ),
    .X(_18601_));
 sky130_fd_sc_hd__a2111o_2 _21282_ (.A1(_18595_),
    .A2(\irq_pending[2] ),
    .B1(_18597_),
    .C1(_18599_),
    .D1(_18601_),
    .X(_18602_));
 sky130_vsdinv _21283_ (.A(\irq_mask[17] ),
    .Y(_18603_));
 sky130_vsdinv _21284_ (.A(\irq_pending[16] ),
    .Y(_18604_));
 sky130_fd_sc_hd__nor2_4 _21285_ (.A(\irq_mask[16] ),
    .B(_18604_),
    .Y(_18605_));
 sky130_vsdinv _21286_ (.A(\irq_mask[19] ),
    .Y(_18606_));
 sky130_fd_sc_hd__and2_1 _21287_ (.A(_18606_),
    .B(\irq_pending[19] ),
    .X(_18607_));
 sky130_vsdinv _21288_ (.A(\irq_mask[18] ),
    .Y(_18608_));
 sky130_fd_sc_hd__and2_1 _21289_ (.A(_18608_),
    .B(\irq_pending[18] ),
    .X(_18609_));
 sky130_fd_sc_hd__a2111o_1 _21290_ (.A1(_18603_),
    .A2(\irq_pending[17] ),
    .B1(_18605_),
    .C1(_18607_),
    .D1(_18609_),
    .X(_18610_));
 sky130_fd_sc_hd__and2b_1 _21291_ (.A_N(\irq_mask[27] ),
    .B(\irq_pending[27] ),
    .X(_18611_));
 sky130_fd_sc_hd__and2b_1 _21292_ (.A_N(\irq_mask[26] ),
    .B(\irq_pending[26] ),
    .X(_18612_));
 sky130_vsdinv _21293_ (.A(\irq_mask[25] ),
    .Y(_18613_));
 sky130_vsdinv _21294_ (.A(\irq_mask[24] ),
    .Y(_18614_));
 sky130_fd_sc_hd__a22o_1 _21295_ (.A1(_18613_),
    .A2(\irq_pending[25] ),
    .B1(_18614_),
    .B2(\irq_pending[24] ),
    .X(_18615_));
 sky130_fd_sc_hd__or3_1 _21296_ (.A(_18611_),
    .B(_18612_),
    .C(_18615_),
    .X(_18616_));
 sky130_vsdinv _21297_ (.A(\irq_mask[23] ),
    .Y(_18617_));
 sky130_fd_sc_hd__and2_1 _21298_ (.A(_18617_),
    .B(\irq_pending[23] ),
    .X(_18618_));
 sky130_fd_sc_hd__and2b_2 _21299_ (.A_N(\irq_mask[22] ),
    .B(\irq_pending[22] ),
    .X(_18619_));
 sky130_vsdinv _21300_ (.A(\irq_mask[21] ),
    .Y(_18620_));
 sky130_vsdinv _21301_ (.A(\irq_mask[20] ),
    .Y(_18621_));
 sky130_fd_sc_hd__a22o_1 _21302_ (.A1(_18620_),
    .A2(\irq_pending[21] ),
    .B1(_18621_),
    .B2(\irq_pending[20] ),
    .X(_18622_));
 sky130_fd_sc_hd__or3_1 _21303_ (.A(_18618_),
    .B(_18619_),
    .C(_18622_),
    .X(_18623_));
 sky130_fd_sc_hd__or4_4 _21304_ (.A(_18602_),
    .B(_18610_),
    .C(_18616_),
    .D(_18623_),
    .X(_18624_));
 sky130_fd_sc_hd__and2b_1 _21305_ (.A_N(\irq_mask[11] ),
    .B(\irq_pending[11] ),
    .X(_18625_));
 sky130_fd_sc_hd__and2b_1 _21306_ (.A_N(\irq_mask[10] ),
    .B(\irq_pending[10] ),
    .X(_18626_));
 sky130_vsdinv _21307_ (.A(\irq_mask[9] ),
    .Y(_18627_));
 sky130_vsdinv _21308_ (.A(\irq_mask[8] ),
    .Y(_18628_));
 sky130_fd_sc_hd__a22o_1 _21309_ (.A1(_18627_),
    .A2(\irq_pending[9] ),
    .B1(_18628_),
    .B2(\irq_pending[8] ),
    .X(_18629_));
 sky130_fd_sc_hd__or3_1 _21310_ (.A(_18625_),
    .B(_18626_),
    .C(_18629_),
    .X(_18630_));
 sky130_fd_sc_hd__and2b_1 _21311_ (.A_N(\irq_mask[7] ),
    .B(\irq_pending[7] ),
    .X(_18631_));
 sky130_fd_sc_hd__and2b_1 _21312_ (.A_N(\irq_mask[6] ),
    .B(\irq_pending[6] ),
    .X(_18632_));
 sky130_vsdinv _21313_ (.A(\irq_mask[5] ),
    .Y(_18633_));
 sky130_vsdinv _21314_ (.A(\irq_mask[4] ),
    .Y(_18634_));
 sky130_fd_sc_hd__a22o_1 _21315_ (.A1(_18633_),
    .A2(\irq_pending[5] ),
    .B1(_18634_),
    .B2(\irq_pending[4] ),
    .X(_18635_));
 sky130_fd_sc_hd__or3_1 _21316_ (.A(_18631_),
    .B(_18632_),
    .C(_18635_),
    .X(_18636_));
 sky130_vsdinv _21317_ (.A(\irq_mask[29] ),
    .Y(_18637_));
 sky130_vsdinv _21318_ (.A(\irq_mask[28] ),
    .Y(_18638_));
 sky130_fd_sc_hd__and2_1 _21319_ (.A(_18638_),
    .B(\irq_pending[28] ),
    .X(_18639_));
 sky130_vsdinv _21320_ (.A(\irq_mask[31] ),
    .Y(_18640_));
 sky130_fd_sc_hd__and2_1 _21321_ (.A(_18640_),
    .B(\irq_pending[31] ),
    .X(_18641_));
 sky130_vsdinv _21322_ (.A(\irq_mask[30] ),
    .Y(_18642_));
 sky130_fd_sc_hd__and2_1 _21323_ (.A(_18642_),
    .B(\irq_pending[30] ),
    .X(_18643_));
 sky130_fd_sc_hd__a2111o_1 _21324_ (.A1(_18637_),
    .A2(\irq_pending[29] ),
    .B1(_18639_),
    .C1(_18641_),
    .D1(_18643_),
    .X(_18644_));
 sky130_vsdinv _21325_ (.A(\irq_mask[13] ),
    .Y(_18645_));
 sky130_vsdinv _21326_ (.A(\irq_mask[12] ),
    .Y(_18646_));
 sky130_fd_sc_hd__and2_1 _21327_ (.A(_18646_),
    .B(\irq_pending[12] ),
    .X(_18647_));
 sky130_vsdinv _21328_ (.A(\irq_mask[15] ),
    .Y(_18648_));
 sky130_fd_sc_hd__and2_1 _21329_ (.A(_18648_),
    .B(\irq_pending[15] ),
    .X(_18649_));
 sky130_vsdinv _21330_ (.A(\irq_mask[14] ),
    .Y(_18650_));
 sky130_fd_sc_hd__and2_1 _21331_ (.A(_18650_),
    .B(\irq_pending[14] ),
    .X(_18651_));
 sky130_fd_sc_hd__a2111o_1 _21332_ (.A1(_18645_),
    .A2(\irq_pending[13] ),
    .B1(_18647_),
    .C1(_18649_),
    .D1(_18651_),
    .X(_18652_));
 sky130_fd_sc_hd__or4_4 _21333_ (.A(_18630_),
    .B(_18636_),
    .C(_18644_),
    .D(_18652_),
    .X(_18653_));
 sky130_fd_sc_hd__nor2_2 _21334_ (.A(_18624_),
    .B(_18653_),
    .Y(_18654_));
 sky130_fd_sc_hd__or4_4 _21335_ (.A(irq_active),
    .B(irq_delay),
    .C(_18594_),
    .D(_18654_),
    .X(_18655_));
 sky130_fd_sc_hd__nor2_2 _21336_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .Y(_18656_));
 sky130_fd_sc_hd__nand2_1 _21337_ (.A(_18655_),
    .B(_18656_),
    .Y(_18657_));
 sky130_vsdinv _21338_ (.A(_18657_),
    .Y(_18658_));
 sky130_vsdinv _21339_ (.A(instr_waitirq),
    .Y(_18659_));
 sky130_fd_sc_hd__nor2_2 _21340_ (.A(_18592_),
    .B(do_waitirq),
    .Y(_18660_));
 sky130_fd_sc_hd__nor2_4 _21341_ (.A(_18659_),
    .B(_18660_),
    .Y(_00309_));
 sky130_vsdinv _21342_ (.A(_00309_),
    .Y(_18661_));
 sky130_fd_sc_hd__nand2_2 _21343_ (.A(_18658_),
    .B(_18661_),
    .Y(_18662_));
 sky130_fd_sc_hd__or2_4 _21344_ (.A(_18593_),
    .B(_18662_),
    .X(_18663_));
 sky130_vsdinv _21345_ (.A(_18663_),
    .Y(_18664_));
 sky130_vsdinv _21346_ (.A(irq_active),
    .Y(_18665_));
 sky130_fd_sc_hd__nand2_1 _21347_ (.A(_18664_),
    .B(_18665_),
    .Y(_18666_));
 sky130_fd_sc_hd__o211a_1 _21348_ (.A1(irq_delay),
    .A2(_18664_),
    .B1(_18549_),
    .C1(_18666_),
    .X(_04065_));
 sky130_vsdinv _21349_ (.A(net330),
    .Y(_18667_));
 sky130_vsdinv _21350_ (.A(net291),
    .Y(_18668_));
 sky130_fd_sc_hd__or4_1 _21351_ (.A(net293),
    .B(net292),
    .C(net279),
    .D(_18668_),
    .X(_18669_));
 sky130_fd_sc_hd__nor3b_4 _21352_ (.A(net302),
    .B(net299),
    .C_N(net300),
    .Y(_18670_));
 sky130_fd_sc_hd__and3b_1 _21353_ (.A_N(net296),
    .B(net285),
    .C(net274),
    .X(_18671_));
 sky130_fd_sc_hd__and4b_1 _21354_ (.A_N(_18669_),
    .B(net301),
    .C(_18670_),
    .D(_18671_),
    .X(_18672_));
 sky130_fd_sc_hd__nand2_4 _21355_ (.A(net101),
    .B(net370),
    .Y(_18673_));
 sky130_fd_sc_hd__or4_4 _21356_ (.A(net298),
    .B(net297),
    .C(net295),
    .D(net294),
    .X(_18674_));
 sky130_fd_sc_hd__nor2_4 _21357_ (.A(_18673_),
    .B(_18674_),
    .Y(_18675_));
 sky130_vsdinv _21358_ (.A(\pcpi_mul.active[0] ),
    .Y(_18676_));
 sky130_vsdinv _21359_ (.A(\pcpi_mul.active[1] ),
    .Y(_18677_));
 sky130_fd_sc_hd__and3_2 _21360_ (.A(_18675_),
    .B(_18676_),
    .C(_18677_),
    .X(_18678_));
 sky130_fd_sc_hd__nand2_4 _21361_ (.A(_18672_),
    .B(_18678_),
    .Y(_18679_));
 sky130_fd_sc_hd__clkbuf_4 _21362_ (.A(_18679_),
    .X(_18680_));
 sky130_fd_sc_hd__nor2_2 _21363_ (.A(_18667_),
    .B(_18680_),
    .Y(_18681_));
 sky130_fd_sc_hd__nor2_1 _21364_ (.A(net278),
    .B(net277),
    .Y(_18682_));
 sky130_vsdinv _21365_ (.A(_18682_),
    .Y(_18683_));
 sky130_fd_sc_hd__nand2_1 _21366_ (.A(net278),
    .B(net277),
    .Y(_18684_));
 sky130_fd_sc_hd__buf_6 _21367_ (.A(\pcpi_mul.rs1[32] ),
    .X(_18685_));
 sky130_fd_sc_hd__buf_6 _21368_ (.A(_18685_),
    .X(_18686_));
 sky130_fd_sc_hd__buf_6 _21369_ (.A(_18686_),
    .X(_18687_));
 sky130_fd_sc_hd__buf_2 _21370_ (.A(_18687_),
    .X(_18688_));
 sky130_fd_sc_hd__buf_2 _21371_ (.A(_18680_),
    .X(_18689_));
 sky130_fd_sc_hd__a32o_1 _21372_ (.A1(_18681_),
    .A2(_18683_),
    .A3(_18684_),
    .B1(_18688_),
    .B2(_18689_),
    .X(_04064_));
 sky130_vsdinv _21373_ (.A(net362),
    .Y(_18690_));
 sky130_fd_sc_hd__nor2_2 _21374_ (.A(_18690_),
    .B(_18680_),
    .Y(_18691_));
 sky130_vsdinv _21375_ (.A(net278),
    .Y(_18692_));
 sky130_fd_sc_hd__buf_6 _21376_ (.A(\pcpi_mul.rs2[32] ),
    .X(_18693_));
 sky130_fd_sc_hd__clkbuf_8 _21377_ (.A(_18693_),
    .X(_18694_));
 sky130_fd_sc_hd__clkbuf_2 _21378_ (.A(_18694_),
    .X(_18695_));
 sky130_fd_sc_hd__clkbuf_2 _21379_ (.A(_18695_),
    .X(_18696_));
 sky130_fd_sc_hd__a32o_1 _21380_ (.A1(_18691_),
    .A2(_18692_),
    .A3(net277),
    .B1(_18696_),
    .B2(_18689_),
    .X(_04063_));
 sky130_fd_sc_hd__buf_2 _21381_ (.A(\cpu_state[4] ),
    .X(_18697_));
 sky130_vsdinv _21382_ (.A(_00333_),
    .Y(_18698_));
 sky130_fd_sc_hd__clkbuf_4 _21383_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_18699_));
 sky130_vsdinv _21384_ (.A(_18699_),
    .Y(_18700_));
 sky130_fd_sc_hd__nor2_2 _21385_ (.A(alu_wait),
    .B(_18700_),
    .Y(_18701_));
 sky130_fd_sc_hd__nor2_1 _21386_ (.A(_18698_),
    .B(_18701_),
    .Y(_18702_));
 sky130_fd_sc_hd__clkbuf_4 _21387_ (.A(_18548_),
    .X(_18703_));
 sky130_fd_sc_hd__o221a_1 _21388_ (.A1(_18697_),
    .A2(_18698_),
    .B1(latched_stalu),
    .B2(_18702_),
    .C1(_18703_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_4 _21389_ (.A(\cpu_state[2] ),
    .X(_18704_));
 sky130_vsdinv _21390_ (.A(_18704_),
    .Y(_18705_));
 sky130_fd_sc_hd__buf_2 _21391_ (.A(_18705_),
    .X(_18706_));
 sky130_fd_sc_hd__buf_2 _21392_ (.A(_18706_),
    .X(_18707_));
 sky130_fd_sc_hd__or4_4 _21393_ (.A(instr_rdinstrh),
    .B(instr_rdinstr),
    .C(instr_rdcycleh),
    .D(instr_rdcycle),
    .X(_18708_));
 sky130_fd_sc_hd__nor2_4 _21394_ (.A(instr_setq),
    .B(instr_getq),
    .Y(_18709_));
 sky130_fd_sc_hd__nand2_2 _21395_ (.A(_18709_),
    .B(_18551_),
    .Y(_18710_));
 sky130_vsdinv _21396_ (.A(_18710_),
    .Y(_18711_));
 sky130_vsdinv _21397_ (.A(instr_timer),
    .Y(_18712_));
 sky130_fd_sc_hd__clkbuf_4 _21398_ (.A(instr_maskirq),
    .X(_18713_));
 sky130_vsdinv _21399_ (.A(_18713_),
    .Y(_18714_));
 sky130_fd_sc_hd__and3_4 _21400_ (.A(_18711_),
    .B(_18712_),
    .C(_18714_),
    .X(_01717_));
 sky130_fd_sc_hd__and2b_1 _21401_ (.A_N(_18708_),
    .B(_01717_),
    .X(_18715_));
 sky130_vsdinv _21402_ (.A(_18715_),
    .Y(_18716_));
 sky130_fd_sc_hd__nor2_1 _21403_ (.A(_18707_),
    .B(_18716_),
    .Y(_18717_));
 sky130_fd_sc_hd__buf_2 _21404_ (.A(\cpu_state[3] ),
    .X(_18718_));
 sky130_fd_sc_hd__nor2_8 _21405_ (.A(\cpu_state[4] ),
    .B(net518),
    .Y(_18719_));
 sky130_fd_sc_hd__clkinv_8 _21406_ (.A(_18719_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _21407_ (.A(_18718_),
    .B(_02542_),
    .Y(_00354_));
 sky130_vsdinv _21408_ (.A(\cpu_state[1] ),
    .Y(_18720_));
 sky130_fd_sc_hd__clkbuf_2 _21409_ (.A(_18720_),
    .X(_18721_));
 sky130_fd_sc_hd__clkbuf_2 _21410_ (.A(_18536_),
    .X(_18722_));
 sky130_fd_sc_hd__a32o_1 _21411_ (.A1(_00354_),
    .A2(_18721_),
    .A3(_18722_),
    .B1(\cpu_state[4] ),
    .B2(alu_wait),
    .X(_18723_));
 sky130_vsdinv _21412_ (.A(instr_sltiu),
    .Y(_18724_));
 sky130_vsdinv _21413_ (.A(instr_slti),
    .Y(_18725_));
 sky130_fd_sc_hd__nand2_1 _21414_ (.A(_18724_),
    .B(_18725_),
    .Y(_18726_));
 sky130_fd_sc_hd__or4_4 _21415_ (.A(instr_and),
    .B(instr_or),
    .C(instr_xor),
    .D(instr_sltu),
    .X(_18727_));
 sky130_fd_sc_hd__or4_4 _21416_ (.A(instr_bgeu),
    .B(instr_bge),
    .C(_18726_),
    .D(_18727_),
    .X(_18728_));
 sky130_fd_sc_hd__or4_4 _21417_ (.A(instr_maskirq),
    .B(_18708_),
    .C(_18710_),
    .D(_18728_),
    .X(_18729_));
 sky130_fd_sc_hd__or4_4 _21418_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_18730_));
 sky130_vsdinv _21419_ (.A(instr_slt),
    .Y(_18731_));
 sky130_vsdinv _21420_ (.A(instr_sll),
    .Y(_18732_));
 sky130_fd_sc_hd__nand2_1 _21421_ (.A(_18731_),
    .B(_18732_),
    .Y(_18733_));
 sky130_fd_sc_hd__or4_4 _21422_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_addi),
    .X(_18734_));
 sky130_fd_sc_hd__or4_4 _21423_ (.A(instr_sub),
    .B(instr_add),
    .C(_18733_),
    .D(_18734_),
    .X(_18735_));
 sky130_fd_sc_hd__or4_4 _21424_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_18736_));
 sky130_fd_sc_hd__nor2_8 _21425_ (.A(instr_auipc),
    .B(instr_lui),
    .Y(_18737_));
 sky130_fd_sc_hd__inv_2 _21426_ (.A(instr_jal),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _21427_ (.A(_18737_),
    .B(_00323_),
    .Y(_00005_));
 sky130_fd_sc_hd__or4_4 _21428_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_18738_));
 sky130_fd_sc_hd__or4_4 _21429_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_18739_));
 sky130_fd_sc_hd__or4_4 _21430_ (.A(instr_sra),
    .B(instr_srl),
    .C(instr_srai),
    .D(instr_srli),
    .X(_18740_));
 sky130_fd_sc_hd__or4_4 _21431_ (.A(_00005_),
    .B(_18738_),
    .C(_18739_),
    .D(_18740_),
    .X(_18741_));
 sky130_fd_sc_hd__or4_4 _21432_ (.A(_18730_),
    .B(_18735_),
    .C(_18736_),
    .D(_18741_),
    .X(_18742_));
 sky130_fd_sc_hd__nor2_4 _21433_ (.A(_18729_),
    .B(_18742_),
    .Y(_00310_));
 sky130_vsdinv _21434_ (.A(net517),
    .Y(_18743_));
 sky130_fd_sc_hd__a21o_1 _21435_ (.A1(_00310_),
    .A2(\pcpi_mul.active[1] ),
    .B1(_18743_),
    .X(_18744_));
 sky130_fd_sc_hd__or3b_1 _21436_ (.A(_18717_),
    .B(_18723_),
    .C_N(_18744_),
    .X(_18745_));
 sky130_vsdinv _21437_ (.A(net511),
    .Y(_18746_));
 sky130_fd_sc_hd__nand2_1 _21438_ (.A(_18745_),
    .B(_18746_),
    .Y(_18747_));
 sky130_fd_sc_hd__o211a_1 _21439_ (.A1(_21142_),
    .A2(_18745_),
    .B1(_18549_),
    .C1(_18747_),
    .X(_04061_));
 sky130_fd_sc_hd__buf_4 _21440_ (.A(\irq_state[0] ),
    .X(_18748_));
 sky130_vsdinv _21441_ (.A(_18748_),
    .Y(_18749_));
 sky130_fd_sc_hd__or2_1 _21442_ (.A(\irq_state[1] ),
    .B(_18720_),
    .X(_18750_));
 sky130_fd_sc_hd__or2_1 _21443_ (.A(_18749_),
    .B(_18750_),
    .X(_18751_));
 sky130_fd_sc_hd__buf_2 _21444_ (.A(_18721_),
    .X(_18752_));
 sky130_fd_sc_hd__buf_1 _21445_ (.A(\irq_state[1] ),
    .X(_18753_));
 sky130_fd_sc_hd__clkbuf_4 _21446_ (.A(_18753_),
    .X(_18754_));
 sky130_fd_sc_hd__nand2_1 _21447_ (.A(_18752_),
    .B(_18754_),
    .Y(_18755_));
 sky130_fd_sc_hd__clkbuf_4 _21448_ (.A(_18533_),
    .X(_18756_));
 sky130_fd_sc_hd__clkbuf_2 _21449_ (.A(_18756_),
    .X(_18757_));
 sky130_fd_sc_hd__clkbuf_4 _21450_ (.A(_18757_),
    .X(_18758_));
 sky130_fd_sc_hd__a21oi_1 _21451_ (.A1(_18751_),
    .A2(_18755_),
    .B1(_18758_),
    .Y(_04060_));
 sky130_fd_sc_hd__buf_1 _21452_ (.A(\irq_state[1] ),
    .X(_18759_));
 sky130_fd_sc_hd__or4_4 _21453_ (.A(_18759_),
    .B(_18748_),
    .C(_18721_),
    .D(_18655_),
    .X(_18760_));
 sky130_fd_sc_hd__clkbuf_4 _21454_ (.A(\irq_state[0] ),
    .X(_18761_));
 sky130_fd_sc_hd__clkbuf_4 _21455_ (.A(_18761_),
    .X(_18762_));
 sky130_fd_sc_hd__nand2_1 _21456_ (.A(_18752_),
    .B(_18762_),
    .Y(_18763_));
 sky130_fd_sc_hd__a21oi_1 _21457_ (.A1(_18760_),
    .A2(_18763_),
    .B1(_18758_),
    .Y(_04059_));
 sky130_vsdinv _21458_ (.A(_00310_),
    .Y(_18764_));
 sky130_fd_sc_hd__nand2_1 _21459_ (.A(_18764_),
    .B(is_lb_lh_lw_lbu_lhu),
    .Y(_18765_));
 sky130_fd_sc_hd__and3_1 _21460_ (.A(_18719_),
    .B(_18721_),
    .C(_18743_),
    .X(_18766_));
 sky130_vsdinv _21461_ (.A(\cpu_state[4] ),
    .Y(_18767_));
 sky130_fd_sc_hd__nor2_2 _21462_ (.A(alu_wait),
    .B(_18767_),
    .Y(_18768_));
 sky130_fd_sc_hd__a21oi_1 _21463_ (.A1(is_sb_sh_sw),
    .A2(_18764_),
    .B1(_18744_),
    .Y(_18769_));
 sky130_fd_sc_hd__a2111oi_2 _21464_ (.A1(_18704_),
    .A2(_18765_),
    .B1(_18766_),
    .C1(_18768_),
    .D1(_18769_),
    .Y(_18770_));
 sky130_vsdinv _21465_ (.A(_18770_),
    .Y(_18771_));
 sky130_vsdinv _21466_ (.A(_18530_),
    .Y(_18772_));
 sky130_fd_sc_hd__nor2_4 _21467_ (.A(_18557_),
    .B(_18772_),
    .Y(_18773_));
 sky130_fd_sc_hd__buf_2 _21468_ (.A(\cpu_state[1] ),
    .X(_18774_));
 sky130_fd_sc_hd__nor2_1 _21469_ (.A(_18774_),
    .B(net518),
    .Y(_00315_));
 sky130_vsdinv _21470_ (.A(_00315_),
    .Y(_18775_));
 sky130_fd_sc_hd__or3_1 _21471_ (.A(\cpu_state[0] ),
    .B(_18718_),
    .C(_18775_),
    .X(_18776_));
 sky130_fd_sc_hd__nor2_8 _21472_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .Y(_00297_));
 sky130_vsdinv _21473_ (.A(_00297_),
    .Y(_18777_));
 sky130_fd_sc_hd__nand2_1 _21474_ (.A(_18701_),
    .B(_18540_),
    .Y(_18778_));
 sky130_fd_sc_hd__or3_2 _21475_ (.A(_00343_),
    .B(_18777_),
    .C(_18778_),
    .X(_18779_));
 sky130_fd_sc_hd__nor2_1 _21476_ (.A(_18776_),
    .B(_18779_),
    .Y(_18780_));
 sky130_fd_sc_hd__and3b_1 _21477_ (.A_N(_00356_),
    .B(_18770_),
    .C(_18773_),
    .X(_18781_));
 sky130_fd_sc_hd__a311o_1 _21478_ (.A1(mem_do_rinst),
    .A2(_18771_),
    .A3(_18773_),
    .B1(_18780_),
    .C1(_18781_),
    .X(_04058_));
 sky130_fd_sc_hd__inv_2 _21479_ (.A(instr_jalr),
    .Y(_02063_));
 sky130_fd_sc_hd__buf_2 _21480_ (.A(instr_jal),
    .X(_18782_));
 sky130_fd_sc_hd__a211o_1 _21481_ (.A1(_18551_),
    .A2(_02063_),
    .B1(_18782_),
    .C1(_18593_),
    .X(_18783_));
 sky130_fd_sc_hd__nor2_1 _21482_ (.A(_18782_),
    .B(_18663_),
    .Y(_18784_));
 sky130_fd_sc_hd__o221a_1 _21483_ (.A1(_18662_),
    .A2(_18783_),
    .B1(mem_do_prefetch),
    .B2(_18784_),
    .C1(_18773_),
    .X(_04057_));
 sky130_fd_sc_hd__nor2_1 _21484_ (.A(net491),
    .B(net478),
    .Y(_18785_));
 sky130_fd_sc_hd__nor2_1 _21485_ (.A(net502),
    .B(net498),
    .Y(_18786_));
 sky130_fd_sc_hd__and3_1 _21486_ (.A(_18785_),
    .B(_18786_),
    .C(_00368_),
    .X(_18787_));
 sky130_fd_sc_hd__buf_4 _21487_ (.A(_18787_),
    .X(_18788_));
 sky130_fd_sc_hd__nor2_8 _21488_ (.A(_01207_),
    .B(_18788_),
    .Y(\cpuregs_rs1[31] ));
 sky130_fd_sc_hd__nor2_1 _21489_ (.A(_18714_),
    .B(_18706_),
    .Y(_18789_));
 sky130_fd_sc_hd__clkbuf_2 _21490_ (.A(_18789_),
    .X(_18790_));
 sky130_fd_sc_hd__clkbuf_2 _21491_ (.A(_18790_),
    .X(_18791_));
 sky130_fd_sc_hd__buf_2 _21492_ (.A(_18791_),
    .X(_18792_));
 sky130_fd_sc_hd__buf_2 _21493_ (.A(_18756_),
    .X(_18793_));
 sky130_fd_sc_hd__buf_4 _21494_ (.A(_18793_),
    .X(_18794_));
 sky130_fd_sc_hd__clkbuf_2 _21495_ (.A(_18790_),
    .X(_18795_));
 sky130_fd_sc_hd__nor2_1 _21496_ (.A(_18640_),
    .B(_18795_),
    .Y(_18796_));
 sky130_fd_sc_hd__a211o_1 _21497_ (.A1(\cpuregs_rs1[31] ),
    .A2(_18792_),
    .B1(_18794_),
    .C1(_18796_),
    .X(_04056_));
 sky130_vsdinv _21498_ (.A(_18789_),
    .Y(_18797_));
 sky130_fd_sc_hd__clkbuf_2 _21499_ (.A(_18797_),
    .X(_18798_));
 sky130_fd_sc_hd__buf_6 _21500_ (.A(_18787_),
    .X(_18799_));
 sky130_fd_sc_hd__nor2_4 _21501_ (.A(_18799_),
    .B(_18797_),
    .Y(_18800_));
 sky130_fd_sc_hd__clkbuf_2 _21502_ (.A(_18800_),
    .X(_18801_));
 sky130_vsdinv _21503_ (.A(_01180_),
    .Y(_18802_));
 sky130_fd_sc_hd__buf_2 _21504_ (.A(_18557_),
    .X(_18803_));
 sky130_fd_sc_hd__buf_2 _21505_ (.A(_18803_),
    .X(_18804_));
 sky130_fd_sc_hd__a221o_1 _21506_ (.A1(\irq_mask[30] ),
    .A2(_18798_),
    .B1(_18801_),
    .B2(_18802_),
    .C1(_18804_),
    .X(_04055_));
 sky130_fd_sc_hd__nor2_8 _21507_ (.A(_01180_),
    .B(net439),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__buf_4 _21508_ (.A(_18799_),
    .X(_18805_));
 sky130_fd_sc_hd__nor2_8 _21509_ (.A(_01153_),
    .B(net434),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__nor2_1 _21510_ (.A(_18637_),
    .B(_18795_),
    .Y(_18806_));
 sky130_fd_sc_hd__a211o_1 _21511_ (.A1(\cpuregs_rs1[29] ),
    .A2(_18792_),
    .B1(_18794_),
    .C1(_18806_),
    .X(_04054_));
 sky130_vsdinv _21512_ (.A(_01126_),
    .Y(_18807_));
 sky130_fd_sc_hd__a221o_1 _21513_ (.A1(\irq_mask[28] ),
    .A2(_18798_),
    .B1(_18801_),
    .B2(_18807_),
    .C1(_18804_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_8 _21514_ (.A(_01126_),
    .B(net439),
    .Y(\cpuregs_rs1[28] ));
 sky130_vsdinv _21515_ (.A(_01099_),
    .Y(_18808_));
 sky130_fd_sc_hd__clkbuf_2 _21516_ (.A(_18803_),
    .X(_18809_));
 sky130_fd_sc_hd__a221o_1 _21517_ (.A1(\irq_mask[27] ),
    .A2(_18798_),
    .B1(_18801_),
    .B2(_18808_),
    .C1(_18809_),
    .X(_04052_));
 sky130_fd_sc_hd__nor2_8 _21518_ (.A(_01099_),
    .B(_18805_),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__buf_6 _21519_ (.A(_18799_),
    .X(_18810_));
 sky130_fd_sc_hd__nor2_8 _21520_ (.A(_01072_),
    .B(_18810_),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__clkbuf_2 _21521_ (.A(_18803_),
    .X(_18811_));
 sky130_fd_sc_hd__clkbuf_2 _21522_ (.A(_18797_),
    .X(_18812_));
 sky130_fd_sc_hd__and2_1 _21523_ (.A(_18812_),
    .B(\irq_mask[26] ),
    .X(_18813_));
 sky130_fd_sc_hd__a211o_1 _21524_ (.A1(\cpuregs_rs1[26] ),
    .A2(_18792_),
    .B1(_18811_),
    .C1(_18813_),
    .X(_04051_));
 sky130_fd_sc_hd__nor2_8 _21525_ (.A(_01045_),
    .B(net433),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__clkbuf_2 _21526_ (.A(_18790_),
    .X(_18814_));
 sky130_fd_sc_hd__nor2_1 _21527_ (.A(_18613_),
    .B(_18814_),
    .Y(_18815_));
 sky130_fd_sc_hd__a211o_1 _21528_ (.A1(\cpuregs_rs1[25] ),
    .A2(_18792_),
    .B1(_18811_),
    .C1(_18815_),
    .X(_04050_));
 sky130_fd_sc_hd__buf_4 _21529_ (.A(_18787_),
    .X(_18816_));
 sky130_fd_sc_hd__nor2_8 _21530_ (.A(_01018_),
    .B(net438),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__nor2_1 _21531_ (.A(_18614_),
    .B(_18814_),
    .Y(_18817_));
 sky130_fd_sc_hd__a211o_1 _21532_ (.A1(\cpuregs_rs1[24] ),
    .A2(_18792_),
    .B1(_18811_),
    .C1(_18817_),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_8 _21533_ (.A(_00991_),
    .B(net433),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__nor2_1 _21534_ (.A(_18617_),
    .B(_18814_),
    .Y(_18818_));
 sky130_fd_sc_hd__a211o_1 _21535_ (.A1(\cpuregs_rs1[23] ),
    .A2(_18792_),
    .B1(_18811_),
    .C1(_18818_),
    .X(_04048_));
 sky130_vsdinv _21536_ (.A(_00964_),
    .Y(_18819_));
 sky130_fd_sc_hd__a221o_1 _21537_ (.A1(\irq_mask[22] ),
    .A2(_18798_),
    .B1(_18801_),
    .B2(_18819_),
    .C1(_18809_),
    .X(_04047_));
 sky130_fd_sc_hd__nor2_8 _21538_ (.A(_00964_),
    .B(net434),
    .Y(\cpuregs_rs1[22] ));
 sky130_vsdinv _21539_ (.A(_00937_),
    .Y(_18820_));
 sky130_fd_sc_hd__a221o_1 _21540_ (.A1(\irq_mask[21] ),
    .A2(_18798_),
    .B1(_18801_),
    .B2(_18820_),
    .C1(_18809_),
    .X(_04046_));
 sky130_fd_sc_hd__nor2_8 _21541_ (.A(_00937_),
    .B(net434),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__nor2_8 _21542_ (.A(_00910_),
    .B(net433),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__buf_2 _21543_ (.A(_18790_),
    .X(_18821_));
 sky130_fd_sc_hd__nor2_1 _21544_ (.A(_18621_),
    .B(_18814_),
    .Y(_18822_));
 sky130_fd_sc_hd__a211o_1 _21545_ (.A1(\cpuregs_rs1[20] ),
    .A2(_18821_),
    .B1(_18811_),
    .C1(_18822_),
    .X(_04045_));
 sky130_vsdinv _21546_ (.A(_00883_),
    .Y(_18823_));
 sky130_fd_sc_hd__a221o_1 _21547_ (.A1(\irq_mask[19] ),
    .A2(_18812_),
    .B1(_18801_),
    .B2(_18823_),
    .C1(_18809_),
    .X(_04044_));
 sky130_fd_sc_hd__nor2_8 _21548_ (.A(_00883_),
    .B(net439),
    .Y(\cpuregs_rs1[19] ));
 sky130_vsdinv _21549_ (.A(_00856_),
    .Y(_18824_));
 sky130_fd_sc_hd__a221o_1 _21550_ (.A1(\irq_mask[18] ),
    .A2(_18812_),
    .B1(_18800_),
    .B2(_18824_),
    .C1(_18809_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_8 _21551_ (.A(_00856_),
    .B(net439),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__nor2_8 _21552_ (.A(_00829_),
    .B(_18810_),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__nor2_1 _21553_ (.A(_18603_),
    .B(_18814_),
    .Y(_18825_));
 sky130_fd_sc_hd__a211o_1 _21554_ (.A1(\cpuregs_rs1[17] ),
    .A2(_18821_),
    .B1(_18811_),
    .C1(_18825_),
    .X(_04042_));
 sky130_vsdinv _21555_ (.A(_00802_),
    .Y(_18826_));
 sky130_fd_sc_hd__a221o_1 _21556_ (.A1(\irq_mask[16] ),
    .A2(_18812_),
    .B1(_18800_),
    .B2(_18826_),
    .C1(_18809_),
    .X(_04041_));
 sky130_fd_sc_hd__nor2_8 _21557_ (.A(_00802_),
    .B(net434),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__nor2_8 _21558_ (.A(_00775_),
    .B(_18816_),
    .Y(\cpuregs_rs1[15] ));
 sky130_fd_sc_hd__clkbuf_2 _21559_ (.A(_18803_),
    .X(_18827_));
 sky130_fd_sc_hd__nor2_1 _21560_ (.A(_18648_),
    .B(_18814_),
    .Y(_18828_));
 sky130_fd_sc_hd__a211o_1 _21561_ (.A1(\cpuregs_rs1[15] ),
    .A2(_18821_),
    .B1(_18827_),
    .C1(_18828_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_8 _21562_ (.A(_00748_),
    .B(_18816_),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__clkbuf_2 _21563_ (.A(_18790_),
    .X(_18829_));
 sky130_fd_sc_hd__nor2_1 _21564_ (.A(_18650_),
    .B(_18829_),
    .Y(_18830_));
 sky130_fd_sc_hd__a211o_1 _21565_ (.A1(\cpuregs_rs1[14] ),
    .A2(_18821_),
    .B1(_18827_),
    .C1(_18830_),
    .X(_04039_));
 sky130_fd_sc_hd__nor2_8 _21566_ (.A(_00721_),
    .B(net433),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__nor2_1 _21567_ (.A(_18645_),
    .B(_18829_),
    .Y(_18831_));
 sky130_fd_sc_hd__a211o_1 _21568_ (.A1(\cpuregs_rs1[13] ),
    .A2(_18821_),
    .B1(_18827_),
    .C1(_18831_),
    .X(_04038_));
 sky130_fd_sc_hd__buf_4 _21569_ (.A(_18799_),
    .X(_18832_));
 sky130_fd_sc_hd__nor2_8 _21570_ (.A(_00694_),
    .B(_18832_),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__nor2_1 _21571_ (.A(_18646_),
    .B(_18829_),
    .Y(_18833_));
 sky130_fd_sc_hd__a211o_1 _21572_ (.A1(\cpuregs_rs1[12] ),
    .A2(_18821_),
    .B1(_18827_),
    .C1(_18833_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_8 _21573_ (.A(_00667_),
    .B(net432),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__clkbuf_2 _21574_ (.A(_18790_),
    .X(_18834_));
 sky130_fd_sc_hd__and2_1 _21575_ (.A(_18797_),
    .B(\irq_mask[11] ),
    .X(_18835_));
 sky130_fd_sc_hd__a211o_1 _21576_ (.A1(\cpuregs_rs1[11] ),
    .A2(_18834_),
    .B1(_18827_),
    .C1(_18835_),
    .X(_04036_));
 sky130_fd_sc_hd__nor2_8 _21577_ (.A(_00640_),
    .B(net432),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__and2_1 _21578_ (.A(_18797_),
    .B(\irq_mask[10] ),
    .X(_18836_));
 sky130_fd_sc_hd__a211o_1 _21579_ (.A1(\cpuregs_rs1[10] ),
    .A2(_18834_),
    .B1(_18827_),
    .C1(_18836_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_8 _21580_ (.A(_00613_),
    .B(_18832_),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__clkbuf_2 _21581_ (.A(_18803_),
    .X(_18837_));
 sky130_fd_sc_hd__nor2_1 _21582_ (.A(_18627_),
    .B(_18829_),
    .Y(_18838_));
 sky130_fd_sc_hd__a211o_1 _21583_ (.A1(\cpuregs_rs1[9] ),
    .A2(_18834_),
    .B1(_18837_),
    .C1(_18838_),
    .X(_04034_));
 sky130_fd_sc_hd__nor2_8 _21584_ (.A(_00586_),
    .B(net438),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__nor2_1 _21585_ (.A(_18628_),
    .B(_18829_),
    .Y(_18839_));
 sky130_fd_sc_hd__a211o_1 _21586_ (.A1(\cpuregs_rs1[8] ),
    .A2(_18834_),
    .B1(_18837_),
    .C1(_18839_),
    .X(_04033_));
 sky130_fd_sc_hd__nor2_8 _21587_ (.A(_00559_),
    .B(net438),
    .Y(\cpuregs_rs1[7] ));
 sky130_vsdinv _21588_ (.A(\irq_mask[7] ),
    .Y(_18840_));
 sky130_fd_sc_hd__nor2_1 _21589_ (.A(_18840_),
    .B(_18829_),
    .Y(_18841_));
 sky130_fd_sc_hd__a211o_1 _21590_ (.A1(\cpuregs_rs1[7] ),
    .A2(_18834_),
    .B1(_18837_),
    .C1(_18841_),
    .X(_04032_));
 sky130_vsdinv _21591_ (.A(_00532_),
    .Y(_18842_));
 sky130_fd_sc_hd__buf_4 _21592_ (.A(_18803_),
    .X(_18843_));
 sky130_fd_sc_hd__a221o_1 _21593_ (.A1(\irq_mask[6] ),
    .A2(_18812_),
    .B1(_18800_),
    .B2(_18842_),
    .C1(_18843_),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_8 _21594_ (.A(_00532_),
    .B(_18805_),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__nor2_8 _21595_ (.A(_00505_),
    .B(net432),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__nor2_1 _21596_ (.A(_18633_),
    .B(_18791_),
    .Y(_18844_));
 sky130_fd_sc_hd__a211o_1 _21597_ (.A1(\cpuregs_rs1[5] ),
    .A2(_18834_),
    .B1(_18837_),
    .C1(_18844_),
    .X(_04030_));
 sky130_fd_sc_hd__nor2_8 _21598_ (.A(_00478_),
    .B(net432),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__nor2_1 _21599_ (.A(_18634_),
    .B(_18791_),
    .Y(_18845_));
 sky130_fd_sc_hd__a211o_1 _21600_ (.A1(\cpuregs_rs1[4] ),
    .A2(_18795_),
    .B1(_18837_),
    .C1(_18845_),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_8 _21601_ (.A(_00451_),
    .B(net438),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__nor2_1 _21602_ (.A(_18600_),
    .B(_18791_),
    .Y(_18846_));
 sky130_fd_sc_hd__a211o_1 _21603_ (.A1(\cpuregs_rs1[3] ),
    .A2(_18795_),
    .B1(_18837_),
    .C1(_18846_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_8 _21604_ (.A(_00424_),
    .B(_18788_),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__nor2_1 _21605_ (.A(_18595_),
    .B(_18791_),
    .Y(_18847_));
 sky130_fd_sc_hd__a211o_1 _21606_ (.A1(\cpuregs_rs1[2] ),
    .A2(_18795_),
    .B1(_18804_),
    .C1(_18847_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_8 _21607_ (.A(_00397_),
    .B(_18799_),
    .Y(\cpuregs_rs1[1] ));
 sky130_vsdinv _21608_ (.A(\irq_mask[1] ),
    .Y(_18848_));
 sky130_fd_sc_hd__nor2_1 _21609_ (.A(_18848_),
    .B(_18791_),
    .Y(_18849_));
 sky130_fd_sc_hd__a211o_1 _21610_ (.A1(\cpuregs_rs1[1] ),
    .A2(_18795_),
    .B1(_18804_),
    .C1(_18849_),
    .X(_04026_));
 sky130_vsdinv _21611_ (.A(_18799_),
    .Y(_18850_));
 sky130_fd_sc_hd__nand2_2 _21612_ (.A(_18850_),
    .B(_00370_),
    .Y(_18851_));
 sky130_fd_sc_hd__nor2_1 _21613_ (.A(_18812_),
    .B(_18851_),
    .Y(_18852_));
 sky130_fd_sc_hd__a211o_1 _21614_ (.A1(\irq_mask[0] ),
    .A2(_18798_),
    .B1(_18804_),
    .C1(_18852_),
    .X(_04025_));
 sky130_vsdinv _21615_ (.A(_18851_),
    .Y(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__clkbuf_2 _21616_ (.A(mem_do_wdata),
    .X(_18853_));
 sky130_fd_sc_hd__buf_6 _21617_ (.A(_18561_),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_1 _21618_ (.A(_18853_),
    .B(_00301_),
    .Y(_18854_));
 sky130_fd_sc_hd__nor2_8 _21619_ (.A(_18532_),
    .B(_18560_),
    .Y(_18855_));
 sky130_fd_sc_hd__nand2_4 _21620_ (.A(_18564_),
    .B(_18855_),
    .Y(_00316_));
 sky130_fd_sc_hd__nor2_8 _21621_ (.A(net408),
    .B(_00316_),
    .Y(_18856_));
 sky130_fd_sc_hd__buf_4 _21622_ (.A(_18856_),
    .X(_18857_));
 sky130_fd_sc_hd__mux2_1 _21623_ (.A0(net166),
    .A1(_18854_),
    .S(_18857_),
    .X(_04024_));
 sky130_vsdinv _21624_ (.A(_00328_),
    .Y(_18858_));
 sky130_fd_sc_hd__and3_1 _21625_ (.A(_18858_),
    .B(_00329_),
    .C(_00330_),
    .X(_18859_));
 sky130_vsdinv _21626_ (.A(_18577_),
    .Y(_18860_));
 sky130_fd_sc_hd__a31o_1 _21627_ (.A1(_18579_),
    .A2(_18581_),
    .A3(_18859_),
    .B1(_18860_),
    .X(_18861_));
 sky130_fd_sc_hd__o211a_1 _21628_ (.A1(_18699_),
    .A2(_18578_),
    .B1(_18549_),
    .C1(_18861_),
    .X(_04023_));
 sky130_fd_sc_hd__buf_2 _21629_ (.A(_18576_),
    .X(_18862_));
 sky130_fd_sc_hd__nand2_1 _21630_ (.A(_18862_),
    .B(\mem_rdata_latched[18] ),
    .Y(_18863_));
 sky130_fd_sc_hd__buf_2 _21631_ (.A(_18860_),
    .X(_00337_));
 sky130_fd_sc_hd__a2bb2o_1 _21632_ (.A1_N(_18863_),
    .A2_N(_18587_),
    .B1(\decoded_rs1[3] ),
    .B2(_00337_),
    .X(_04022_));
 sky130_fd_sc_hd__nand2_1 _21633_ (.A(_18862_),
    .B(\mem_rdata_latched[17] ),
    .Y(_18864_));
 sky130_fd_sc_hd__a2bb2o_1 _21634_ (.A1_N(_18864_),
    .A2_N(_18587_),
    .B1(\decoded_rs1[2] ),
    .B2(_00337_),
    .X(_04021_));
 sky130_fd_sc_hd__nand2_1 _21635_ (.A(_18862_),
    .B(\mem_rdata_latched[16] ),
    .Y(_18865_));
 sky130_fd_sc_hd__a2bb2o_1 _21636_ (.A1_N(_18865_),
    .A2_N(_18587_),
    .B1(\decoded_rs1[1] ),
    .B2(_00337_),
    .X(_04020_));
 sky130_fd_sc_hd__nand2_1 _21637_ (.A(_18862_),
    .B(\mem_rdata_latched[15] ),
    .Y(_18866_));
 sky130_fd_sc_hd__a2bb2o_1 _21638_ (.A1_N(_18866_),
    .A2_N(_18587_),
    .B1(\decoded_rs1[0] ),
    .B2(_00337_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_2 _21639_ (.A(_18757_),
    .X(_18867_));
 sky130_fd_sc_hd__nor2_2 _21640_ (.A(decoder_pseudo_trigger),
    .B(_18594_),
    .Y(_18868_));
 sky130_vsdinv _21641_ (.A(_18868_),
    .Y(_18869_));
 sky130_fd_sc_hd__buf_2 _21642_ (.A(_18869_),
    .X(_18870_));
 sky130_fd_sc_hd__clkbuf_4 _21643_ (.A(_18870_),
    .X(_18871_));
 sky130_fd_sc_hd__inv_2 _21644_ (.A(\mem_rdata_q[14] ),
    .Y(_00334_));
 sky130_vsdinv _21645_ (.A(\mem_rdata_q[13] ),
    .Y(_18872_));
 sky130_fd_sc_hd__clkbuf_2 _21646_ (.A(_18872_),
    .X(_18873_));
 sky130_vsdinv _21647_ (.A(\mem_rdata_q[12] ),
    .Y(_18874_));
 sky130_fd_sc_hd__or3_4 _21648_ (.A(_00334_),
    .B(_18873_),
    .C(_18874_),
    .X(_18875_));
 sky130_vsdinv _21649_ (.A(\mem_rdata_q[31] ),
    .Y(_18876_));
 sky130_vsdinv _21650_ (.A(\mem_rdata_q[30] ),
    .Y(_18877_));
 sky130_vsdinv _21651_ (.A(\mem_rdata_q[29] ),
    .Y(_18878_));
 sky130_fd_sc_hd__and3_1 _21652_ (.A(_18876_),
    .B(_18877_),
    .C(_18878_),
    .X(_18879_));
 sky130_vsdinv _21653_ (.A(\mem_rdata_q[27] ),
    .Y(_18880_));
 sky130_vsdinv _21654_ (.A(decoder_pseudo_trigger),
    .Y(_18881_));
 sky130_fd_sc_hd__and3_1 _21655_ (.A(_18880_),
    .B(_18881_),
    .C(_18592_),
    .X(_18882_));
 sky130_fd_sc_hd__nor2_1 _21656_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .Y(_18883_));
 sky130_vsdinv _21657_ (.A(\mem_rdata_q[25] ),
    .Y(_18884_));
 sky130_fd_sc_hd__and2_1 _21658_ (.A(_18883_),
    .B(_18884_),
    .X(_18885_));
 sky130_fd_sc_hd__and3_1 _21659_ (.A(_18879_),
    .B(_18882_),
    .C(_18885_),
    .X(_18886_));
 sky130_fd_sc_hd__nand2_2 _21660_ (.A(_18886_),
    .B(is_alu_reg_reg),
    .Y(_18887_));
 sky130_fd_sc_hd__o2bb2a_1 _21661_ (.A1_N(instr_and),
    .A2_N(_18871_),
    .B1(_18875_),
    .B2(_18887_),
    .X(_18888_));
 sky130_fd_sc_hd__nor2_1 _21662_ (.A(_18867_),
    .B(_18888_),
    .Y(_04018_));
 sky130_fd_sc_hd__buf_2 _21663_ (.A(\mem_rdata_q[12] ),
    .X(_18889_));
 sky130_fd_sc_hd__or3_4 _21664_ (.A(_18889_),
    .B(_00334_),
    .C(_18873_),
    .X(_18890_));
 sky130_fd_sc_hd__o2bb2a_1 _21665_ (.A1_N(instr_or),
    .A2_N(_18871_),
    .B1(_18890_),
    .B2(_18887_),
    .X(_18891_));
 sky130_fd_sc_hd__nor2_1 _21666_ (.A(_18867_),
    .B(_18891_),
    .Y(_04017_));
 sky130_vsdinv _21667_ (.A(is_alu_reg_reg),
    .Y(_18892_));
 sky130_fd_sc_hd__buf_2 _21668_ (.A(\mem_rdata_q[14] ),
    .X(_18893_));
 sky130_fd_sc_hd__and3_1 _21669_ (.A(_18873_),
    .B(_18893_),
    .C(\mem_rdata_q[12] ),
    .X(_18894_));
 sky130_vsdinv _21670_ (.A(_18894_),
    .Y(_18895_));
 sky130_fd_sc_hd__and3_1 _21671_ (.A(_18878_),
    .B(_18881_),
    .C(_18592_),
    .X(_18896_));
 sky130_vsdinv _21672_ (.A(_18896_),
    .Y(_18897_));
 sky130_fd_sc_hd__buf_2 _21673_ (.A(\mem_rdata_q[25] ),
    .X(_18898_));
 sky130_fd_sc_hd__nand2_1 _21674_ (.A(_18883_),
    .B(_18880_),
    .Y(_18899_));
 sky130_fd_sc_hd__or4_4 _21675_ (.A(\mem_rdata_q[31] ),
    .B(_18877_),
    .C(_18898_),
    .D(_18899_),
    .X(_18900_));
 sky130_fd_sc_hd__nor2_1 _21676_ (.A(_18897_),
    .B(_18900_),
    .Y(_18901_));
 sky130_vsdinv _21677_ (.A(_18901_),
    .Y(_18902_));
 sky130_fd_sc_hd__or3_1 _21678_ (.A(_18892_),
    .B(_18895_),
    .C(_18902_),
    .X(_18903_));
 sky130_fd_sc_hd__clkbuf_2 _21679_ (.A(_18870_),
    .X(_18904_));
 sky130_fd_sc_hd__clkbuf_4 _21680_ (.A(_18904_),
    .X(_18905_));
 sky130_fd_sc_hd__nand2_1 _21681_ (.A(_18905_),
    .B(instr_sra),
    .Y(_18906_));
 sky130_fd_sc_hd__a21oi_1 _21682_ (.A1(_18903_),
    .A2(_18906_),
    .B1(_18758_),
    .Y(_04016_));
 sky130_fd_sc_hd__clkbuf_2 _21683_ (.A(_18886_),
    .X(_18907_));
 sky130_fd_sc_hd__buf_2 _21684_ (.A(_18870_),
    .X(_18908_));
 sky130_fd_sc_hd__a32o_1 _21685_ (.A1(_18907_),
    .A2(is_alu_reg_reg),
    .A3(_18894_),
    .B1(instr_srl),
    .B2(_18908_),
    .X(_18909_));
 sky130_fd_sc_hd__and2_1 _21686_ (.A(_18909_),
    .B(_18703_),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_2 _21687_ (.A(_18870_),
    .X(_18910_));
 sky130_fd_sc_hd__and3_1 _21688_ (.A(_18873_),
    .B(_18874_),
    .C(_18893_),
    .X(_18911_));
 sky130_vsdinv _21689_ (.A(_18911_),
    .Y(_18912_));
 sky130_fd_sc_hd__o2bb2a_1 _21690_ (.A1_N(instr_xor),
    .A2_N(_18910_),
    .B1(_18912_),
    .B2(_18887_),
    .X(_18913_));
 sky130_fd_sc_hd__nor2_1 _21691_ (.A(_18867_),
    .B(_18913_),
    .Y(_04014_));
 sky130_fd_sc_hd__nor2_1 _21692_ (.A(\mem_rdata_q[14] ),
    .B(_18872_),
    .Y(_18914_));
 sky130_fd_sc_hd__nand2_1 _21693_ (.A(_18914_),
    .B(_18889_),
    .Y(_18915_));
 sky130_fd_sc_hd__o2bb2a_1 _21694_ (.A1_N(instr_sltu),
    .A2_N(_18910_),
    .B1(_18915_),
    .B2(_18887_),
    .X(_18916_));
 sky130_fd_sc_hd__nor2_1 _21695_ (.A(_18867_),
    .B(_18916_),
    .Y(_04013_));
 sky130_fd_sc_hd__clkbuf_2 _21696_ (.A(_18868_),
    .X(_18917_));
 sky130_fd_sc_hd__clkbuf_2 _21697_ (.A(_18917_),
    .X(_18918_));
 sky130_fd_sc_hd__nand2_2 _21698_ (.A(_18914_),
    .B(_18874_),
    .Y(_18919_));
 sky130_fd_sc_hd__o22a_1 _21699_ (.A1(_18731_),
    .A2(_18918_),
    .B1(_18919_),
    .B2(_18887_),
    .X(_18920_));
 sky130_fd_sc_hd__nor2_1 _21700_ (.A(_18867_),
    .B(_18920_),
    .Y(_04012_));
 sky130_fd_sc_hd__clkbuf_2 _21701_ (.A(_18757_),
    .X(_18921_));
 sky130_fd_sc_hd__clkbuf_2 _21702_ (.A(_18917_),
    .X(_18922_));
 sky130_fd_sc_hd__and3_1 _21703_ (.A(_00334_),
    .B(_18873_),
    .C(\mem_rdata_q[12] ),
    .X(_18923_));
 sky130_vsdinv _21704_ (.A(_18923_),
    .Y(_18924_));
 sky130_fd_sc_hd__o22a_1 _21705_ (.A1(_18732_),
    .A2(_18922_),
    .B1(_18924_),
    .B2(_18887_),
    .X(_18925_));
 sky130_fd_sc_hd__nor2_1 _21706_ (.A(_18921_),
    .B(_18925_),
    .Y(_04011_));
 sky130_fd_sc_hd__and3_2 _21707_ (.A(_00334_),
    .B(_18872_),
    .C(_18874_),
    .X(_18926_));
 sky130_vsdinv _21708_ (.A(_18926_),
    .Y(_18927_));
 sky130_fd_sc_hd__or3_2 _21709_ (.A(_18892_),
    .B(_18927_),
    .C(_18902_),
    .X(_18928_));
 sky130_fd_sc_hd__nand2_1 _21710_ (.A(_18905_),
    .B(instr_sub),
    .Y(_18929_));
 sky130_fd_sc_hd__a21oi_1 _21711_ (.A1(_18928_),
    .A2(_18929_),
    .B1(_18758_),
    .Y(_04010_));
 sky130_fd_sc_hd__buf_2 _21712_ (.A(_18870_),
    .X(_18930_));
 sky130_fd_sc_hd__a32o_1 _21713_ (.A1(_18907_),
    .A2(is_alu_reg_reg),
    .A3(_18926_),
    .B1(instr_add),
    .B2(_18930_),
    .X(_18931_));
 sky130_fd_sc_hd__and2_1 _21714_ (.A(_18931_),
    .B(_18543_),
    .X(_04009_));
 sky130_vsdinv _21715_ (.A(is_alu_reg_imm),
    .Y(_18932_));
 sky130_fd_sc_hd__nor2_4 _21716_ (.A(_18932_),
    .B(_18869_),
    .Y(_18933_));
 sky130_vsdinv _21717_ (.A(_18933_),
    .Y(_18934_));
 sky130_fd_sc_hd__o2bb2a_1 _21718_ (.A1_N(instr_andi),
    .A2_N(_18910_),
    .B1(_18875_),
    .B2(_18934_),
    .X(_18935_));
 sky130_fd_sc_hd__nor2_1 _21719_ (.A(_18921_),
    .B(_18935_),
    .Y(_04008_));
 sky130_fd_sc_hd__o2bb2a_1 _21720_ (.A1_N(instr_ori),
    .A2_N(_18910_),
    .B1(_18890_),
    .B2(_18934_),
    .X(_18936_));
 sky130_fd_sc_hd__nor2_1 _21721_ (.A(_18921_),
    .B(_18936_),
    .Y(_04007_));
 sky130_fd_sc_hd__a22o_1 _21722_ (.A1(instr_xori),
    .A2(_18930_),
    .B1(_18933_),
    .B2(_18911_),
    .X(_18937_));
 sky130_fd_sc_hd__and2_1 _21723_ (.A(_18937_),
    .B(_18543_),
    .X(_04006_));
 sky130_fd_sc_hd__o22a_1 _21724_ (.A1(_18724_),
    .A2(_18922_),
    .B1(_18915_),
    .B2(_18934_),
    .X(_18938_));
 sky130_fd_sc_hd__nor2_1 _21725_ (.A(_18921_),
    .B(_18938_),
    .Y(_04005_));
 sky130_fd_sc_hd__o22a_1 _21726_ (.A1(_18725_),
    .A2(_18922_),
    .B1(_18919_),
    .B2(_18934_),
    .X(_18939_));
 sky130_fd_sc_hd__nor2_1 _21727_ (.A(_18921_),
    .B(_18939_),
    .Y(_04004_));
 sky130_fd_sc_hd__a22o_1 _21728_ (.A1(instr_addi),
    .A2(_18930_),
    .B1(_18933_),
    .B2(_18926_),
    .X(_18940_));
 sky130_fd_sc_hd__and2_1 _21729_ (.A(_18940_),
    .B(_18543_),
    .X(_04003_));
 sky130_vsdinv _21730_ (.A(instr_bgeu),
    .Y(_18941_));
 sky130_fd_sc_hd__nand2_2 _21731_ (.A(_18917_),
    .B(_18699_),
    .Y(_18942_));
 sky130_fd_sc_hd__o22a_1 _21732_ (.A1(_18941_),
    .A2(_18922_),
    .B1(_18942_),
    .B2(_18875_),
    .X(_18943_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(_18921_),
    .B(_18943_),
    .Y(_04002_));
 sky130_fd_sc_hd__clkbuf_2 _21734_ (.A(_18757_),
    .X(_18944_));
 sky130_fd_sc_hd__o2bb2a_1 _21735_ (.A1_N(instr_bltu),
    .A2_N(_18910_),
    .B1(_18942_),
    .B2(_18890_),
    .X(_18945_));
 sky130_fd_sc_hd__nor2_1 _21736_ (.A(_18944_),
    .B(_18945_),
    .Y(_04001_));
 sky130_fd_sc_hd__o2bb2a_1 _21737_ (.A1_N(instr_bge),
    .A2_N(_18910_),
    .B1(_18942_),
    .B2(_18895_),
    .X(_18946_));
 sky130_fd_sc_hd__nor2_1 _21738_ (.A(_18944_),
    .B(_18946_),
    .Y(_04000_));
 sky130_fd_sc_hd__o2bb2a_1 _21739_ (.A1_N(instr_blt),
    .A2_N(_18908_),
    .B1(_18942_),
    .B2(_18912_),
    .X(_18947_));
 sky130_fd_sc_hd__nor2_1 _21740_ (.A(_18944_),
    .B(_18947_),
    .Y(_03999_));
 sky130_vsdinv _21741_ (.A(instr_bne),
    .Y(_18948_));
 sky130_fd_sc_hd__o22a_1 _21742_ (.A1(_18948_),
    .A2(_18922_),
    .B1(_18942_),
    .B2(_18924_),
    .X(_18949_));
 sky130_fd_sc_hd__nor2_1 _21743_ (.A(_18944_),
    .B(_18949_),
    .Y(_03998_));
 sky130_fd_sc_hd__o2bb2a_1 _21744_ (.A1_N(instr_beq),
    .A2_N(_18908_),
    .B1(_18942_),
    .B2(_18927_),
    .X(_18950_));
 sky130_fd_sc_hd__nor2_1 _21745_ (.A(_18944_),
    .B(_18950_),
    .Y(_03997_));
 sky130_vsdinv _21746_ (.A(\pcpi_timeout_counter[3] ),
    .Y(_18951_));
 sky130_fd_sc_hd__nor2_1 _21747_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .Y(_18952_));
 sky130_vsdinv _21748_ (.A(_18952_),
    .Y(_18953_));
 sky130_fd_sc_hd__nor2_2 _21749_ (.A(\pcpi_timeout_counter[2] ),
    .B(_18953_),
    .Y(_18954_));
 sky130_fd_sc_hd__o21bai_1 _21750_ (.A1(_18951_),
    .A2(_18954_),
    .B1_N(_18673_),
    .Y(_03996_));
 sky130_fd_sc_hd__a21o_1 _21751_ (.A1(_18953_),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_18673_),
    .X(_18955_));
 sky130_fd_sc_hd__a21o_1 _21752_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(_18954_),
    .B1(_18955_),
    .X(_03995_));
 sky130_fd_sc_hd__o21a_1 _21753_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_18952_),
    .X(_18956_));
 sky130_fd_sc_hd__a211o_1 _21754_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_18673_),
    .C1(_18956_),
    .X(_03994_));
 sky130_fd_sc_hd__nand2_1 _21755_ (.A(_18954_),
    .B(_18951_),
    .Y(_18957_));
 sky130_vsdinv _21756_ (.A(\pcpi_timeout_counter[0] ),
    .Y(_18958_));
 sky130_fd_sc_hd__a21o_1 _21757_ (.A1(_18957_),
    .A2(_18958_),
    .B1(_18673_),
    .X(_03993_));
 sky130_fd_sc_hd__nor2_4 _21758_ (.A(_18704_),
    .B(_18718_),
    .Y(_18959_));
 sky130_fd_sc_hd__buf_2 _21759_ (.A(_18722_),
    .X(_18960_));
 sky130_fd_sc_hd__and3_4 _21760_ (.A(_18959_),
    .B(_18767_),
    .C(_18960_),
    .X(_01706_));
 sky130_fd_sc_hd__buf_4 _21761_ (.A(_18721_),
    .X(_18961_));
 sky130_vsdinv _21762_ (.A(\cpu_state[0] ),
    .Y(_18962_));
 sky130_fd_sc_hd__and3_1 _21763_ (.A(_00291_),
    .B(_18961_),
    .C(_18962_),
    .X(_18963_));
 sky130_fd_sc_hd__a32o_1 _21764_ (.A1(_18534_),
    .A2(_01706_),
    .A3(_18963_),
    .B1(_18773_),
    .B2(_18853_),
    .X(_03992_));
 sky130_vsdinv _21765_ (.A(mem_do_prefetch),
    .Y(_18964_));
 sky130_fd_sc_hd__nor2_4 _21766_ (.A(_18964_),
    .B(_18573_),
    .Y(_00296_));
 sky130_vsdinv _21767_ (.A(_00296_),
    .Y(_18965_));
 sky130_fd_sc_hd__and3_1 _21768_ (.A(_18535_),
    .B(_18541_),
    .C(\cpu_state[6] ),
    .X(_18966_));
 sky130_fd_sc_hd__a22o_1 _21769_ (.A1(mem_do_rdata),
    .A2(_18773_),
    .B1(_18965_),
    .B2(_18966_),
    .X(_03991_));
 sky130_fd_sc_hd__buf_2 _21770_ (.A(_18752_),
    .X(_18967_));
 sky130_fd_sc_hd__clkbuf_2 _21771_ (.A(_18774_),
    .X(_18968_));
 sky130_fd_sc_hd__or2_1 _21772_ (.A(\reg_next_pc[31] ),
    .B(_18968_),
    .X(_18969_));
 sky130_fd_sc_hd__o211a_1 _21773_ (.A1(_02530_),
    .A2(_18967_),
    .B1(_18549_),
    .C1(_18969_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_4 _21774_ (.A(_18752_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_2 _21775_ (.A(_18548_),
    .X(_18970_));
 sky130_fd_sc_hd__clkbuf_4 _21776_ (.A(_18774_),
    .X(_18971_));
 sky130_fd_sc_hd__clkbuf_2 _21777_ (.A(_18971_),
    .X(_18972_));
 sky130_fd_sc_hd__or2_1 _21778_ (.A(_18972_),
    .B(\reg_next_pc[30] ),
    .X(_18973_));
 sky130_fd_sc_hd__o211a_1 _21779_ (.A1(_00322_),
    .A2(_02529_),
    .B1(_18970_),
    .C1(_18973_),
    .X(_03989_));
 sky130_fd_sc_hd__or2_1 _21780_ (.A(_18972_),
    .B(\reg_next_pc[29] ),
    .X(_18974_));
 sky130_fd_sc_hd__o211a_1 _21781_ (.A1(_00322_),
    .A2(_02527_),
    .B1(_18970_),
    .C1(_18974_),
    .X(_03988_));
 sky130_fd_sc_hd__or2_1 _21782_ (.A(_18972_),
    .B(\reg_next_pc[28] ),
    .X(_18975_));
 sky130_fd_sc_hd__o211a_1 _21783_ (.A1(_00322_),
    .A2(_02526_),
    .B1(_18970_),
    .C1(_18975_),
    .X(_03987_));
 sky130_fd_sc_hd__or2_1 _21784_ (.A(_18972_),
    .B(\reg_next_pc[27] ),
    .X(_18976_));
 sky130_fd_sc_hd__o211a_1 _21785_ (.A1(_00322_),
    .A2(_02525_),
    .B1(_18970_),
    .C1(_18976_),
    .X(_03986_));
 sky130_fd_sc_hd__or2_1 _21786_ (.A(_18972_),
    .B(\reg_next_pc[26] ),
    .X(_18977_));
 sky130_fd_sc_hd__o211a_1 _21787_ (.A1(_00322_),
    .A2(_02524_),
    .B1(_18970_),
    .C1(_18977_),
    .X(_03985_));
 sky130_fd_sc_hd__buf_2 _21788_ (.A(_18961_),
    .X(_18978_));
 sky130_fd_sc_hd__or2_1 _21789_ (.A(_18972_),
    .B(\reg_next_pc[25] ),
    .X(_18979_));
 sky130_fd_sc_hd__o211a_1 _21790_ (.A1(_18978_),
    .A2(_02523_),
    .B1(_18970_),
    .C1(_18979_),
    .X(_03984_));
 sky130_fd_sc_hd__clkbuf_4 _21791_ (.A(_18547_),
    .X(_18980_));
 sky130_fd_sc_hd__clkbuf_2 _21792_ (.A(_18980_),
    .X(_18981_));
 sky130_fd_sc_hd__buf_1 _21793_ (.A(_18971_),
    .X(_18982_));
 sky130_fd_sc_hd__or2_1 _21794_ (.A(_18982_),
    .B(\reg_next_pc[24] ),
    .X(_18983_));
 sky130_fd_sc_hd__o211a_1 _21795_ (.A1(_18978_),
    .A2(_02522_),
    .B1(_18981_),
    .C1(_18983_),
    .X(_03983_));
 sky130_fd_sc_hd__or2_1 _21796_ (.A(_18982_),
    .B(\reg_next_pc[23] ),
    .X(_18984_));
 sky130_fd_sc_hd__o211a_1 _21797_ (.A1(_18978_),
    .A2(_02521_),
    .B1(_18981_),
    .C1(_18984_),
    .X(_03982_));
 sky130_fd_sc_hd__or2_1 _21798_ (.A(_18982_),
    .B(\reg_next_pc[22] ),
    .X(_18985_));
 sky130_fd_sc_hd__o211a_1 _21799_ (.A1(_18978_),
    .A2(_02520_),
    .B1(_18981_),
    .C1(_18985_),
    .X(_03981_));
 sky130_fd_sc_hd__or2_1 _21800_ (.A(_18982_),
    .B(\reg_next_pc[21] ),
    .X(_18986_));
 sky130_fd_sc_hd__o211a_1 _21801_ (.A1(_18978_),
    .A2(_02519_),
    .B1(_18981_),
    .C1(_18986_),
    .X(_03980_));
 sky130_fd_sc_hd__or2_1 _21802_ (.A(_18982_),
    .B(\reg_next_pc[20] ),
    .X(_18987_));
 sky130_fd_sc_hd__o211a_1 _21803_ (.A1(_18978_),
    .A2(_02518_),
    .B1(_18981_),
    .C1(_18987_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_4 _21804_ (.A(_18961_),
    .X(_18988_));
 sky130_fd_sc_hd__or2_1 _21805_ (.A(_18982_),
    .B(\reg_next_pc[19] ),
    .X(_18989_));
 sky130_fd_sc_hd__o211a_1 _21806_ (.A1(_18988_),
    .A2(_02516_),
    .B1(_18981_),
    .C1(_18989_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_4 _21807_ (.A(_18980_),
    .X(_18990_));
 sky130_fd_sc_hd__buf_2 _21808_ (.A(_18774_),
    .X(_18991_));
 sky130_fd_sc_hd__or2_1 _21809_ (.A(_18991_),
    .B(\reg_next_pc[18] ),
    .X(_18992_));
 sky130_fd_sc_hd__o211a_1 _21810_ (.A1(_18988_),
    .A2(_02515_),
    .B1(_18990_),
    .C1(_18992_),
    .X(_03977_));
 sky130_fd_sc_hd__or2_1 _21811_ (.A(_18991_),
    .B(\reg_next_pc[17] ),
    .X(_18993_));
 sky130_fd_sc_hd__o211a_1 _21812_ (.A1(_18988_),
    .A2(_02514_),
    .B1(_18990_),
    .C1(_18993_),
    .X(_03976_));
 sky130_fd_sc_hd__or2_1 _21813_ (.A(_18991_),
    .B(\reg_next_pc[16] ),
    .X(_18994_));
 sky130_fd_sc_hd__o211a_1 _21814_ (.A1(_18988_),
    .A2(_02513_),
    .B1(_18990_),
    .C1(_18994_),
    .X(_03975_));
 sky130_fd_sc_hd__or2_1 _21815_ (.A(_18991_),
    .B(\reg_next_pc[15] ),
    .X(_18995_));
 sky130_fd_sc_hd__o211a_1 _21816_ (.A1(_18988_),
    .A2(_02512_),
    .B1(_18990_),
    .C1(_18995_),
    .X(_03974_));
 sky130_fd_sc_hd__or2_1 _21817_ (.A(_18991_),
    .B(\reg_next_pc[14] ),
    .X(_18996_));
 sky130_fd_sc_hd__o211a_1 _21818_ (.A1(_18988_),
    .A2(_02511_),
    .B1(_18990_),
    .C1(_18996_),
    .X(_03973_));
 sky130_fd_sc_hd__buf_2 _21819_ (.A(_18961_),
    .X(_18997_));
 sky130_fd_sc_hd__or2_1 _21820_ (.A(_18991_),
    .B(\reg_next_pc[13] ),
    .X(_18998_));
 sky130_fd_sc_hd__o211a_1 _21821_ (.A1(_18997_),
    .A2(_02510_),
    .B1(_18990_),
    .C1(_18998_),
    .X(_03972_));
 sky130_fd_sc_hd__clkbuf_2 _21822_ (.A(_18980_),
    .X(_18999_));
 sky130_fd_sc_hd__clkbuf_2 _21823_ (.A(_18774_),
    .X(_19000_));
 sky130_fd_sc_hd__or2_1 _21824_ (.A(_19000_),
    .B(\reg_next_pc[12] ),
    .X(_19001_));
 sky130_fd_sc_hd__o211a_1 _21825_ (.A1(_18997_),
    .A2(_02509_),
    .B1(_18999_),
    .C1(_19001_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_1 _21826_ (.A(_19000_),
    .B(\reg_next_pc[11] ),
    .X(_19002_));
 sky130_fd_sc_hd__o211a_1 _21827_ (.A1(_18997_),
    .A2(_02508_),
    .B1(_18999_),
    .C1(_19002_),
    .X(_03970_));
 sky130_fd_sc_hd__or2_1 _21828_ (.A(_19000_),
    .B(\reg_next_pc[10] ),
    .X(_19003_));
 sky130_fd_sc_hd__o211a_1 _21829_ (.A1(_18997_),
    .A2(_02507_),
    .B1(_18999_),
    .C1(_19003_),
    .X(_03969_));
 sky130_fd_sc_hd__or2_1 _21830_ (.A(_19000_),
    .B(\reg_next_pc[9] ),
    .X(_19004_));
 sky130_fd_sc_hd__o211a_1 _21831_ (.A1(_18997_),
    .A2(_02537_),
    .B1(_18999_),
    .C1(_19004_),
    .X(_03968_));
 sky130_fd_sc_hd__or2_1 _21832_ (.A(_19000_),
    .B(\reg_next_pc[8] ),
    .X(_19005_));
 sky130_fd_sc_hd__o211a_1 _21833_ (.A1(_18997_),
    .A2(_02536_),
    .B1(_18999_),
    .C1(_19005_),
    .X(_03967_));
 sky130_fd_sc_hd__buf_2 _21834_ (.A(_18961_),
    .X(_19006_));
 sky130_fd_sc_hd__or2_1 _21835_ (.A(_19000_),
    .B(\reg_next_pc[7] ),
    .X(_19007_));
 sky130_fd_sc_hd__o211a_1 _21836_ (.A1(_19006_),
    .A2(_02535_),
    .B1(_18999_),
    .C1(_19007_),
    .X(_03966_));
 sky130_fd_sc_hd__buf_2 _21837_ (.A(_18980_),
    .X(_19008_));
 sky130_fd_sc_hd__or2_1 _21838_ (.A(_18968_),
    .B(\reg_next_pc[6] ),
    .X(_19009_));
 sky130_fd_sc_hd__o211a_1 _21839_ (.A1(_19006_),
    .A2(_02534_),
    .B1(_19008_),
    .C1(_19009_),
    .X(_03965_));
 sky130_fd_sc_hd__or2_1 _21840_ (.A(_18968_),
    .B(\reg_next_pc[5] ),
    .X(_19010_));
 sky130_fd_sc_hd__o211a_1 _21841_ (.A1(_19006_),
    .A2(_02533_),
    .B1(_19008_),
    .C1(_19010_),
    .X(_03964_));
 sky130_fd_sc_hd__inv_2 _21842_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _21843_ (.A(_18967_),
    .B(_01471_),
    .Y(_19011_));
 sky130_fd_sc_hd__o211a_1 _21844_ (.A1(_19006_),
    .A2(_02532_),
    .B1(_19008_),
    .C1(_19011_),
    .X(_03963_));
 sky130_fd_sc_hd__or2_1 _21845_ (.A(_18968_),
    .B(\reg_next_pc[3] ),
    .X(_19012_));
 sky130_fd_sc_hd__o211a_1 _21846_ (.A1(_19006_),
    .A2(_02531_),
    .B1(_19008_),
    .C1(_19012_),
    .X(_03962_));
 sky130_fd_sc_hd__or2_1 _21847_ (.A(_18968_),
    .B(\reg_next_pc[2] ),
    .X(_19013_));
 sky130_fd_sc_hd__o211a_1 _21848_ (.A1(_19006_),
    .A2(_02528_),
    .B1(_19008_),
    .C1(_19013_),
    .X(_03961_));
 sky130_fd_sc_hd__or2_1 _21849_ (.A(_18968_),
    .B(\reg_next_pc[1] ),
    .X(_19014_));
 sky130_fd_sc_hd__o211a_1 _21850_ (.A1(_18967_),
    .A2(_02517_),
    .B1(_19008_),
    .C1(_19014_),
    .X(_03960_));
 sky130_fd_sc_hd__clkbuf_4 _21851_ (.A(_18774_),
    .X(_19015_));
 sky130_fd_sc_hd__clkbuf_4 _21852_ (.A(_19015_),
    .X(_19016_));
 sky130_fd_sc_hd__buf_2 _21853_ (.A(_18980_),
    .X(_19017_));
 sky130_vsdinv _21854_ (.A(_02581_),
    .Y(_19018_));
 sky130_fd_sc_hd__clkbuf_4 _21855_ (.A(_18971_),
    .X(_19019_));
 sky130_fd_sc_hd__nand2_1 _21856_ (.A(_19018_),
    .B(_19019_),
    .Y(_19020_));
 sky130_fd_sc_hd__o211a_1 _21857_ (.A1(_19016_),
    .A2(\reg_pc[31] ),
    .B1(_19017_),
    .C1(_19020_),
    .X(_03959_));
 sky130_vsdinv _21858_ (.A(_02580_),
    .Y(_19021_));
 sky130_fd_sc_hd__nand2_1 _21859_ (.A(_19021_),
    .B(_19019_),
    .Y(_19022_));
 sky130_fd_sc_hd__o211a_1 _21860_ (.A1(_19016_),
    .A2(\reg_pc[30] ),
    .B1(_19017_),
    .C1(_19022_),
    .X(_03958_));
 sky130_vsdinv _21861_ (.A(_02579_),
    .Y(_19023_));
 sky130_fd_sc_hd__nand2_1 _21862_ (.A(_19023_),
    .B(_19019_),
    .Y(_19024_));
 sky130_fd_sc_hd__o211a_1 _21863_ (.A1(_19016_),
    .A2(\reg_pc[29] ),
    .B1(_19017_),
    .C1(_19024_),
    .X(_03957_));
 sky130_vsdinv _21864_ (.A(_02578_),
    .Y(_19025_));
 sky130_fd_sc_hd__nand2_1 _21865_ (.A(_19025_),
    .B(_19019_),
    .Y(_19026_));
 sky130_fd_sc_hd__o211a_1 _21866_ (.A1(_19016_),
    .A2(\reg_pc[28] ),
    .B1(_19017_),
    .C1(_19026_),
    .X(_03956_));
 sky130_vsdinv _21867_ (.A(_02577_),
    .Y(_19027_));
 sky130_fd_sc_hd__nand2_1 _21868_ (.A(_19027_),
    .B(_19019_),
    .Y(_19028_));
 sky130_fd_sc_hd__o211a_1 _21869_ (.A1(_19016_),
    .A2(\reg_pc[27] ),
    .B1(_19017_),
    .C1(_19028_),
    .X(_03955_));
 sky130_fd_sc_hd__clkbuf_2 _21870_ (.A(_19015_),
    .X(_19029_));
 sky130_vsdinv _21871_ (.A(_02576_),
    .Y(_19030_));
 sky130_fd_sc_hd__clkbuf_2 _21872_ (.A(_19015_),
    .X(_19031_));
 sky130_fd_sc_hd__nand2_1 _21873_ (.A(_19030_),
    .B(_19031_),
    .Y(_19032_));
 sky130_fd_sc_hd__o211a_1 _21874_ (.A1(_19029_),
    .A2(\reg_pc[26] ),
    .B1(_19017_),
    .C1(_19032_),
    .X(_03954_));
 sky130_fd_sc_hd__clkbuf_2 _21875_ (.A(_18980_),
    .X(_19033_));
 sky130_vsdinv _21876_ (.A(_02575_),
    .Y(_19034_));
 sky130_fd_sc_hd__nand2_1 _21877_ (.A(_19034_),
    .B(_19031_),
    .Y(_19035_));
 sky130_fd_sc_hd__o211a_1 _21878_ (.A1(_19029_),
    .A2(\reg_pc[25] ),
    .B1(_19033_),
    .C1(_19035_),
    .X(_03953_));
 sky130_vsdinv _21879_ (.A(_02574_),
    .Y(_19036_));
 sky130_fd_sc_hd__nand2_1 _21880_ (.A(_19036_),
    .B(_19031_),
    .Y(_19037_));
 sky130_fd_sc_hd__o211a_1 _21881_ (.A1(_19029_),
    .A2(\reg_pc[24] ),
    .B1(_19033_),
    .C1(_19037_),
    .X(_03952_));
 sky130_vsdinv _21882_ (.A(_02573_),
    .Y(_19038_));
 sky130_fd_sc_hd__nand2_1 _21883_ (.A(_19038_),
    .B(_19031_),
    .Y(_19039_));
 sky130_fd_sc_hd__o211a_1 _21884_ (.A1(_19029_),
    .A2(\reg_pc[23] ),
    .B1(_19033_),
    .C1(_19039_),
    .X(_03951_));
 sky130_vsdinv _21885_ (.A(_02572_),
    .Y(_19040_));
 sky130_fd_sc_hd__nand2_1 _21886_ (.A(_19040_),
    .B(_19031_),
    .Y(_19041_));
 sky130_fd_sc_hd__o211a_1 _21887_ (.A1(_19029_),
    .A2(\reg_pc[22] ),
    .B1(_19033_),
    .C1(_19041_),
    .X(_03950_));
 sky130_vsdinv _21888_ (.A(_02570_),
    .Y(_19042_));
 sky130_fd_sc_hd__nand2_1 _21889_ (.A(_19042_),
    .B(_19031_),
    .Y(_19043_));
 sky130_fd_sc_hd__o211a_1 _21890_ (.A1(_19029_),
    .A2(\reg_pc[21] ),
    .B1(_19033_),
    .C1(_19043_),
    .X(_03949_));
 sky130_fd_sc_hd__clkbuf_2 _21891_ (.A(_19015_),
    .X(_19044_));
 sky130_vsdinv _21892_ (.A(_02569_),
    .Y(_19045_));
 sky130_fd_sc_hd__clkbuf_2 _21893_ (.A(_18971_),
    .X(_19046_));
 sky130_fd_sc_hd__nand2_1 _21894_ (.A(_19045_),
    .B(_19046_),
    .Y(_19047_));
 sky130_fd_sc_hd__o211a_1 _21895_ (.A1(_19044_),
    .A2(\reg_pc[20] ),
    .B1(_19033_),
    .C1(_19047_),
    .X(_03948_));
 sky130_fd_sc_hd__buf_4 _21896_ (.A(_18541_),
    .X(_19048_));
 sky130_fd_sc_hd__clkbuf_4 _21897_ (.A(_19048_),
    .X(_19049_));
 sky130_vsdinv _21898_ (.A(_02568_),
    .Y(_19050_));
 sky130_fd_sc_hd__nand2_1 _21899_ (.A(_19050_),
    .B(_19046_),
    .Y(_19051_));
 sky130_fd_sc_hd__o211a_1 _21900_ (.A1(_19044_),
    .A2(\reg_pc[19] ),
    .B1(_19049_),
    .C1(_19051_),
    .X(_03947_));
 sky130_vsdinv _21901_ (.A(_02567_),
    .Y(_19052_));
 sky130_fd_sc_hd__nand2_1 _21902_ (.A(_19052_),
    .B(_19046_),
    .Y(_19053_));
 sky130_fd_sc_hd__o211a_1 _21903_ (.A1(_19044_),
    .A2(\reg_pc[18] ),
    .B1(_19049_),
    .C1(_19053_),
    .X(_03946_));
 sky130_vsdinv _21904_ (.A(_02566_),
    .Y(_19054_));
 sky130_fd_sc_hd__nand2_1 _21905_ (.A(_19054_),
    .B(_19046_),
    .Y(_19055_));
 sky130_fd_sc_hd__o211a_1 _21906_ (.A1(_19044_),
    .A2(\reg_pc[17] ),
    .B1(_19049_),
    .C1(_19055_),
    .X(_03945_));
 sky130_vsdinv _21907_ (.A(_02565_),
    .Y(_19056_));
 sky130_fd_sc_hd__nand2_1 _21908_ (.A(_19056_),
    .B(_19046_),
    .Y(_19057_));
 sky130_fd_sc_hd__o211a_1 _21909_ (.A1(_19044_),
    .A2(\reg_pc[16] ),
    .B1(_19049_),
    .C1(_19057_),
    .X(_03944_));
 sky130_vsdinv _21910_ (.A(_02564_),
    .Y(_19058_));
 sky130_fd_sc_hd__nand2_1 _21911_ (.A(_19058_),
    .B(_19046_),
    .Y(_19059_));
 sky130_fd_sc_hd__o211a_1 _21912_ (.A1(_19044_),
    .A2(\reg_pc[15] ),
    .B1(_19049_),
    .C1(_19059_),
    .X(_03943_));
 sky130_fd_sc_hd__clkbuf_2 _21913_ (.A(_19015_),
    .X(_19060_));
 sky130_vsdinv _21914_ (.A(_02563_),
    .Y(_19061_));
 sky130_fd_sc_hd__clkbuf_2 _21915_ (.A(_18971_),
    .X(_19062_));
 sky130_fd_sc_hd__nand2_1 _21916_ (.A(_19061_),
    .B(_19062_),
    .Y(_19063_));
 sky130_fd_sc_hd__o211a_1 _21917_ (.A1(_19060_),
    .A2(\reg_pc[14] ),
    .B1(_19049_),
    .C1(_19063_),
    .X(_03942_));
 sky130_fd_sc_hd__clkbuf_2 _21918_ (.A(_19048_),
    .X(_19064_));
 sky130_vsdinv _21919_ (.A(_02562_),
    .Y(_19065_));
 sky130_fd_sc_hd__nand2_1 _21920_ (.A(_19065_),
    .B(_19062_),
    .Y(_19066_));
 sky130_fd_sc_hd__o211a_1 _21921_ (.A1(_19060_),
    .A2(\reg_pc[13] ),
    .B1(_19064_),
    .C1(_19066_),
    .X(_03941_));
 sky130_vsdinv _21922_ (.A(_02561_),
    .Y(_19067_));
 sky130_fd_sc_hd__nand2_1 _21923_ (.A(_19067_),
    .B(_19062_),
    .Y(_19068_));
 sky130_fd_sc_hd__o211a_1 _21924_ (.A1(_19060_),
    .A2(\reg_pc[12] ),
    .B1(_19064_),
    .C1(_19068_),
    .X(_03940_));
 sky130_vsdinv _21925_ (.A(_02589_),
    .Y(_19069_));
 sky130_fd_sc_hd__nand2_1 _21926_ (.A(_19069_),
    .B(_19062_),
    .Y(_19070_));
 sky130_fd_sc_hd__o211a_1 _21927_ (.A1(_19060_),
    .A2(\reg_pc[11] ),
    .B1(_19064_),
    .C1(_19070_),
    .X(_03939_));
 sky130_vsdinv _21928_ (.A(_02588_),
    .Y(_19071_));
 sky130_fd_sc_hd__nand2_1 _21929_ (.A(_19071_),
    .B(_19062_),
    .Y(_19072_));
 sky130_fd_sc_hd__o211a_1 _21930_ (.A1(_19060_),
    .A2(\reg_pc[10] ),
    .B1(_19064_),
    .C1(_19072_),
    .X(_03938_));
 sky130_vsdinv _21931_ (.A(_02587_),
    .Y(_19073_));
 sky130_fd_sc_hd__nand2_1 _21932_ (.A(_19073_),
    .B(_19062_),
    .Y(_19074_));
 sky130_fd_sc_hd__o211a_1 _21933_ (.A1(_19060_),
    .A2(\reg_pc[9] ),
    .B1(_19064_),
    .C1(_19074_),
    .X(_03937_));
 sky130_fd_sc_hd__buf_2 _21934_ (.A(_19015_),
    .X(_19075_));
 sky130_vsdinv _21935_ (.A(_02586_),
    .Y(_19076_));
 sky130_fd_sc_hd__clkbuf_4 _21936_ (.A(_18971_),
    .X(_19077_));
 sky130_fd_sc_hd__nand2_1 _21937_ (.A(_19076_),
    .B(_19077_),
    .Y(_19078_));
 sky130_fd_sc_hd__o211a_1 _21938_ (.A1(_19075_),
    .A2(\reg_pc[8] ),
    .B1(_19064_),
    .C1(_19078_),
    .X(_03936_));
 sky130_fd_sc_hd__clkbuf_2 _21939_ (.A(_19048_),
    .X(_19079_));
 sky130_vsdinv _21940_ (.A(_02585_),
    .Y(_19080_));
 sky130_fd_sc_hd__nand2_1 _21941_ (.A(_19080_),
    .B(_19077_),
    .Y(_19081_));
 sky130_fd_sc_hd__o211a_1 _21942_ (.A1(_19075_),
    .A2(\reg_pc[7] ),
    .B1(_19079_),
    .C1(_19081_),
    .X(_03935_));
 sky130_vsdinv _21943_ (.A(_02584_),
    .Y(_19082_));
 sky130_fd_sc_hd__nand2_1 _21944_ (.A(_19082_),
    .B(_19077_),
    .Y(_19083_));
 sky130_fd_sc_hd__o211a_1 _21945_ (.A1(_19075_),
    .A2(\reg_pc[6] ),
    .B1(_19079_),
    .C1(_19083_),
    .X(_03934_));
 sky130_vsdinv _21946_ (.A(_02583_),
    .Y(_19084_));
 sky130_fd_sc_hd__nand2_1 _21947_ (.A(_19084_),
    .B(_19077_),
    .Y(_19085_));
 sky130_fd_sc_hd__o211a_1 _21948_ (.A1(_19075_),
    .A2(\reg_pc[5] ),
    .B1(_19079_),
    .C1(_19085_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _21949_ (.A(_19019_),
    .B(_01475_),
    .Y(_19086_));
 sky130_fd_sc_hd__o211a_1 _21950_ (.A1(_19075_),
    .A2(\reg_pc[4] ),
    .B1(_19079_),
    .C1(_19086_),
    .X(_03932_));
 sky130_fd_sc_hd__inv_2 _21951_ (.A(_01475_),
    .Y(_02582_));
 sky130_vsdinv _21952_ (.A(\reg_pc[3] ),
    .Y(_19087_));
 sky130_fd_sc_hd__nand2_1 _21953_ (.A(_18752_),
    .B(_19087_),
    .Y(_19088_));
 sky130_fd_sc_hd__o211a_1 _21954_ (.A1(_18967_),
    .A2(_02571_),
    .B1(_19079_),
    .C1(_19088_),
    .X(_03931_));
 sky130_fd_sc_hd__inv_2 _21955_ (.A(_02560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _21956_ (.A(_01561_),
    .B(_19077_),
    .Y(_19089_));
 sky130_fd_sc_hd__o211a_1 _21957_ (.A1(_19075_),
    .A2(\reg_pc[2] ),
    .B1(_19079_),
    .C1(_19089_),
    .X(_03930_));
 sky130_fd_sc_hd__buf_6 _21958_ (.A(_19048_),
    .X(_19090_));
 sky130_vsdinv _21959_ (.A(\reg_pc[1] ),
    .Y(_19091_));
 sky130_fd_sc_hd__nand2_1 _21960_ (.A(_18752_),
    .B(_19091_),
    .Y(_19092_));
 sky130_fd_sc_hd__o211a_1 _21961_ (.A1(_18967_),
    .A2(_02590_),
    .B1(_19090_),
    .C1(_19092_),
    .X(_03929_));
 sky130_fd_sc_hd__nand2_2 _21962_ (.A(\count_instr[36] ),
    .B(\count_instr[35] ),
    .Y(_19093_));
 sky130_fd_sc_hd__and2_1 _21963_ (.A(\count_instr[39] ),
    .B(\count_instr[38] ),
    .X(_19094_));
 sky130_fd_sc_hd__nand2_1 _21964_ (.A(_19094_),
    .B(\count_instr[37] ),
    .Y(_19095_));
 sky130_vsdinv _21965_ (.A(\count_instr[25] ),
    .Y(_19096_));
 sky130_vsdinv _21966_ (.A(\count_instr[16] ),
    .Y(_19097_));
 sky130_vsdinv _21967_ (.A(\count_instr[14] ),
    .Y(_19098_));
 sky130_fd_sc_hd__nand2_1 _21968_ (.A(\count_instr[4] ),
    .B(\count_instr[3] ),
    .Y(_19099_));
 sky130_vsdinv _21969_ (.A(\count_instr[12] ),
    .Y(_19100_));
 sky130_vsdinv _21970_ (.A(\count_instr[11] ),
    .Y(_19101_));
 sky130_vsdinv _21971_ (.A(\count_instr[7] ),
    .Y(_19102_));
 sky130_vsdinv _21972_ (.A(\count_instr[6] ),
    .Y(_19103_));
 sky130_fd_sc_hd__or4_4 _21973_ (.A(_19100_),
    .B(_19101_),
    .C(_19102_),
    .D(_19103_),
    .X(_19104_));
 sky130_vsdinv _21974_ (.A(\count_instr[10] ),
    .Y(_19105_));
 sky130_vsdinv _21975_ (.A(\count_instr[9] ),
    .Y(_19106_));
 sky130_vsdinv _21976_ (.A(\count_instr[8] ),
    .Y(_19107_));
 sky130_vsdinv _21977_ (.A(\count_instr[5] ),
    .Y(_19108_));
 sky130_vsdinv _21978_ (.A(\count_instr[2] ),
    .Y(_19109_));
 sky130_vsdinv _21979_ (.A(\count_instr[1] ),
    .Y(_19110_));
 sky130_vsdinv _21980_ (.A(\count_instr[0] ),
    .Y(_19111_));
 sky130_fd_sc_hd__or4_4 _21981_ (.A(_19108_),
    .B(_19109_),
    .C(_19110_),
    .D(_19111_),
    .X(_19112_));
 sky130_fd_sc_hd__or4_4 _21982_ (.A(_19105_),
    .B(_19106_),
    .C(_19107_),
    .D(_19112_),
    .X(_19113_));
 sky130_fd_sc_hd__nor3_1 _21983_ (.A(_19099_),
    .B(_19104_),
    .C(_19113_),
    .Y(_19114_));
 sky130_vsdinv _21984_ (.A(_19114_),
    .Y(_19115_));
 sky130_fd_sc_hd__or3b_4 _21985_ (.A(_19115_),
    .B(_18663_),
    .C_N(\count_instr[13] ),
    .X(_19116_));
 sky130_fd_sc_hd__nor2_2 _21986_ (.A(_19098_),
    .B(_19116_),
    .Y(_19117_));
 sky130_fd_sc_hd__nand2_1 _21987_ (.A(_19117_),
    .B(\count_instr[15] ),
    .Y(_19118_));
 sky130_fd_sc_hd__nor2_1 _21988_ (.A(_19097_),
    .B(_19118_),
    .Y(_19119_));
 sky130_fd_sc_hd__and3_2 _21989_ (.A(_19119_),
    .B(\count_instr[18] ),
    .C(\count_instr[17] ),
    .X(_19120_));
 sky130_vsdinv _21990_ (.A(\count_instr[20] ),
    .Y(_19121_));
 sky130_vsdinv _21991_ (.A(\count_instr[19] ),
    .Y(_19122_));
 sky130_fd_sc_hd__nor2_2 _21992_ (.A(_19121_),
    .B(_19122_),
    .Y(_19123_));
 sky130_fd_sc_hd__and4_1 _21993_ (.A(\count_instr[24] ),
    .B(\count_instr[23] ),
    .C(\count_instr[22] ),
    .D(\count_instr[21] ),
    .X(_19124_));
 sky130_fd_sc_hd__nand3_4 _21994_ (.A(_19120_),
    .B(_19123_),
    .C(_19124_),
    .Y(_19125_));
 sky130_fd_sc_hd__nor3b_4 _21995_ (.A(_19096_),
    .B(_19125_),
    .C_N(\count_instr[26] ),
    .Y(_19126_));
 sky130_vsdinv _21996_ (.A(\count_instr[27] ),
    .Y(_19127_));
 sky130_vsdinv _21997_ (.A(\count_instr[31] ),
    .Y(_19128_));
 sky130_vsdinv _21998_ (.A(\count_instr[30] ),
    .Y(_19129_));
 sky130_vsdinv _21999_ (.A(\count_instr[29] ),
    .Y(_19130_));
 sky130_vsdinv _22000_ (.A(\count_instr[28] ),
    .Y(_19131_));
 sky130_fd_sc_hd__or4_4 _22001_ (.A(_19128_),
    .B(_19129_),
    .C(_19130_),
    .D(_19131_),
    .X(_19132_));
 sky130_fd_sc_hd__nor2_2 _22002_ (.A(_19127_),
    .B(_19132_),
    .Y(_19133_));
 sky130_fd_sc_hd__and3_1 _22003_ (.A(\count_instr[34] ),
    .B(\count_instr[33] ),
    .C(\count_instr[32] ),
    .X(_19134_));
 sky130_fd_sc_hd__nand3_4 _22004_ (.A(_19126_),
    .B(_19133_),
    .C(_19134_),
    .Y(_19135_));
 sky130_fd_sc_hd__nor3_4 _22005_ (.A(_19093_),
    .B(_19095_),
    .C(_19135_),
    .Y(_19136_));
 sky130_fd_sc_hd__and3_1 _22006_ (.A(\count_instr[42] ),
    .B(\count_instr[41] ),
    .C(\count_instr[40] ),
    .X(_19137_));
 sky130_vsdinv _22007_ (.A(\count_instr[49] ),
    .Y(_19138_));
 sky130_vsdinv _22008_ (.A(\count_instr[48] ),
    .Y(_19139_));
 sky130_vsdinv _22009_ (.A(\count_instr[47] ),
    .Y(_19140_));
 sky130_vsdinv _22010_ (.A(\count_instr[46] ),
    .Y(_19141_));
 sky130_vsdinv _22011_ (.A(\count_instr[45] ),
    .Y(_19142_));
 sky130_vsdinv _22012_ (.A(\count_instr[44] ),
    .Y(_19143_));
 sky130_fd_sc_hd__or4_4 _22013_ (.A(_19140_),
    .B(_19141_),
    .C(_19142_),
    .D(_19143_),
    .X(_19144_));
 sky130_fd_sc_hd__nor3_2 _22014_ (.A(_19138_),
    .B(_19139_),
    .C(_19144_),
    .Y(_19145_));
 sky130_fd_sc_hd__and4_1 _22015_ (.A(_19136_),
    .B(\count_instr[43] ),
    .C(_19137_),
    .D(_19145_),
    .X(_19146_));
 sky130_vsdinv _22016_ (.A(\count_instr[52] ),
    .Y(_19147_));
 sky130_vsdinv _22017_ (.A(\count_instr[51] ),
    .Y(_19148_));
 sky130_fd_sc_hd__nor2_2 _22018_ (.A(_19147_),
    .B(_19148_),
    .Y(_19149_));
 sky130_fd_sc_hd__and3_1 _22019_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .C(\count_instr[53] ),
    .X(_19150_));
 sky130_fd_sc_hd__and4_1 _22020_ (.A(_19146_),
    .B(\count_instr[50] ),
    .C(_19149_),
    .D(_19150_),
    .X(_19151_));
 sky130_fd_sc_hd__clkbuf_2 _22021_ (.A(_19151_),
    .X(_19152_));
 sky130_fd_sc_hd__and3_1 _22022_ (.A(\count_instr[58] ),
    .B(\count_instr[57] ),
    .C(\count_instr[56] ),
    .X(_19153_));
 sky130_vsdinv _22023_ (.A(\count_instr[60] ),
    .Y(_19154_));
 sky130_vsdinv _22024_ (.A(\count_instr[59] ),
    .Y(_19155_));
 sky130_fd_sc_hd__nor2_4 _22025_ (.A(_19154_),
    .B(_19155_),
    .Y(_19156_));
 sky130_fd_sc_hd__and3_1 _22026_ (.A(_19156_),
    .B(\count_instr[63] ),
    .C(\count_instr[62] ),
    .X(_19157_));
 sky130_fd_sc_hd__clkbuf_2 _22027_ (.A(_18756_),
    .X(_19158_));
 sky130_fd_sc_hd__a41o_1 _22028_ (.A1(_19152_),
    .A2(\count_instr[61] ),
    .A3(_19153_),
    .A4(_19157_),
    .B1(_19158_),
    .X(_19159_));
 sky130_vsdinv _22029_ (.A(\count_instr[43] ),
    .Y(_19160_));
 sky130_fd_sc_hd__nor2_2 _22030_ (.A(_19160_),
    .B(_19144_),
    .Y(_19161_));
 sky130_fd_sc_hd__nand3_4 _22031_ (.A(_19136_),
    .B(_19137_),
    .C(_19161_),
    .Y(_19162_));
 sky130_vsdinv _22032_ (.A(\count_instr[50] ),
    .Y(_19163_));
 sky130_fd_sc_hd__nor2_1 _22033_ (.A(_19163_),
    .B(_19138_),
    .Y(_19164_));
 sky130_fd_sc_hd__nor3b_4 _22034_ (.A(_19139_),
    .B(_19162_),
    .C_N(_19164_),
    .Y(_19165_));
 sky130_fd_sc_hd__and4_1 _22035_ (.A(_19165_),
    .B(_19149_),
    .C(_19150_),
    .D(_19153_),
    .X(_19166_));
 sky130_fd_sc_hd__clkbuf_2 _22036_ (.A(_19166_),
    .X(_19167_));
 sky130_vsdinv _22037_ (.A(\count_instr[62] ),
    .Y(_19168_));
 sky130_vsdinv _22038_ (.A(\count_instr[61] ),
    .Y(_19169_));
 sky130_fd_sc_hd__nor2_1 _22039_ (.A(_19168_),
    .B(_19169_),
    .Y(_19170_));
 sky130_fd_sc_hd__a31oi_1 _22040_ (.A1(_19167_),
    .A2(_19156_),
    .A3(_19170_),
    .B1(\count_instr[63] ),
    .Y(_19171_));
 sky130_fd_sc_hd__nor2_1 _22041_ (.A(_19159_),
    .B(_19171_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand3_1 _22042_ (.A(_19167_),
    .B(\count_instr[61] ),
    .C(_19156_),
    .Y(_19172_));
 sky130_fd_sc_hd__a41o_1 _22043_ (.A1(_19152_),
    .A2(_19153_),
    .A3(_19156_),
    .A4(_19170_),
    .B1(_18793_),
    .X(_19173_));
 sky130_fd_sc_hd__a21oi_1 _22044_ (.A1(_19172_),
    .A2(_19168_),
    .B1(_19173_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_1 _22045_ (.A(_19167_),
    .B(_19156_),
    .Y(_19174_));
 sky130_fd_sc_hd__buf_4 _22046_ (.A(_18547_),
    .X(_19175_));
 sky130_fd_sc_hd__nand2_1 _22047_ (.A(_19172_),
    .B(_19175_),
    .Y(_19176_));
 sky130_fd_sc_hd__a21oi_1 _22048_ (.A1(_19169_),
    .A2(_19174_),
    .B1(_19176_),
    .Y(_03926_));
 sky130_fd_sc_hd__and3_1 _22049_ (.A(_19151_),
    .B(\count_instr[59] ),
    .C(_19153_),
    .X(_19177_));
 sky130_fd_sc_hd__a21oi_1 _22050_ (.A1(_19167_),
    .A2(_19156_),
    .B1(_18843_),
    .Y(_19178_));
 sky130_fd_sc_hd__o21a_1 _22051_ (.A1(\count_instr[60] ),
    .A2(_19177_),
    .B1(_19178_),
    .X(_03925_));
 sky130_fd_sc_hd__clkbuf_4 _22052_ (.A(_18757_),
    .X(_19179_));
 sky130_fd_sc_hd__nor2_1 _22053_ (.A(\count_instr[59] ),
    .B(_19167_),
    .Y(_19180_));
 sky130_fd_sc_hd__nor3_1 _22054_ (.A(_19179_),
    .B(_19177_),
    .C(_19180_),
    .Y(_03924_));
 sky130_fd_sc_hd__a31o_1 _22055_ (.A1(_19152_),
    .A2(\count_instr[57] ),
    .A3(\count_instr[56] ),
    .B1(\count_instr[58] ),
    .X(_19181_));
 sky130_fd_sc_hd__nor3b_1 _22056_ (.A(_19179_),
    .B(_19167_),
    .C_N(_19181_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand2_1 _22057_ (.A(_19152_),
    .B(\count_instr[56] ),
    .Y(_19182_));
 sky130_vsdinv _22058_ (.A(\count_instr[57] ),
    .Y(_19183_));
 sky130_fd_sc_hd__a31o_1 _22059_ (.A1(_19152_),
    .A2(\count_instr[57] ),
    .A3(\count_instr[56] ),
    .B1(_19158_),
    .X(_19184_));
 sky130_fd_sc_hd__a21oi_1 _22060_ (.A1(_19182_),
    .A2(_19183_),
    .B1(_19184_),
    .Y(_03922_));
 sky130_vsdinv _22061_ (.A(_19152_),
    .Y(_19185_));
 sky130_vsdinv _22062_ (.A(\count_instr[56] ),
    .Y(_19186_));
 sky130_fd_sc_hd__nand2_1 _22063_ (.A(_19185_),
    .B(_19186_),
    .Y(_19187_));
 sky130_fd_sc_hd__clkbuf_2 _22064_ (.A(_18541_),
    .X(_19188_));
 sky130_fd_sc_hd__buf_2 _22065_ (.A(_19188_),
    .X(_19189_));
 sky130_fd_sc_hd__and3_1 _22066_ (.A(_19187_),
    .B(_19189_),
    .C(_19182_),
    .X(_03921_));
 sky130_fd_sc_hd__and3_1 _22067_ (.A(_19146_),
    .B(\count_instr[50] ),
    .C(_19149_),
    .X(_19190_));
 sky130_fd_sc_hd__nand3_1 _22068_ (.A(_19190_),
    .B(\count_instr[54] ),
    .C(\count_instr[53] ),
    .Y(_19191_));
 sky130_vsdinv _22069_ (.A(\count_instr[55] ),
    .Y(_19192_));
 sky130_fd_sc_hd__nand2_1 _22070_ (.A(_19191_),
    .B(_19192_),
    .Y(_19193_));
 sky130_fd_sc_hd__and3_1 _22071_ (.A(_19193_),
    .B(_19189_),
    .C(_19185_),
    .X(_03920_));
 sky130_fd_sc_hd__a31o_1 _22072_ (.A1(_19165_),
    .A2(\count_instr[53] ),
    .A3(_19149_),
    .B1(\count_instr[54] ),
    .X(_19194_));
 sky130_fd_sc_hd__clkbuf_4 _22073_ (.A(_18542_),
    .X(_19195_));
 sky130_fd_sc_hd__and3_1 _22074_ (.A(_19194_),
    .B(_19191_),
    .C(_19195_),
    .X(_03919_));
 sky130_vsdinv _22075_ (.A(_19190_),
    .Y(_19196_));
 sky130_vsdinv _22076_ (.A(\count_instr[53] ),
    .Y(_19197_));
 sky130_fd_sc_hd__nand2_1 _22077_ (.A(_19196_),
    .B(_19197_),
    .Y(_19198_));
 sky130_fd_sc_hd__nand2_1 _22078_ (.A(_19190_),
    .B(\count_instr[53] ),
    .Y(_19199_));
 sky130_fd_sc_hd__and3_1 _22079_ (.A(_19198_),
    .B(_19189_),
    .C(_19199_),
    .X(_03918_));
 sky130_vsdinv _22080_ (.A(_19165_),
    .Y(_19200_));
 sky130_fd_sc_hd__nor2_1 _22081_ (.A(_19148_),
    .B(_19200_),
    .Y(_19201_));
 sky130_fd_sc_hd__o211a_1 _22082_ (.A1(\count_instr[52] ),
    .A2(_19201_),
    .B1(_19090_),
    .C1(_19196_),
    .X(_03917_));
 sky130_fd_sc_hd__nor2_1 _22083_ (.A(_18843_),
    .B(_19201_),
    .Y(_19202_));
 sky130_fd_sc_hd__o21a_1 _22084_ (.A1(\count_instr[51] ),
    .A2(_19165_),
    .B1(_19202_),
    .X(_03916_));
 sky130_vsdinv _22085_ (.A(_19146_),
    .Y(_19203_));
 sky130_fd_sc_hd__nand2_1 _22086_ (.A(_19203_),
    .B(_19163_),
    .Y(_19204_));
 sky130_fd_sc_hd__and3_1 _22087_ (.A(_19200_),
    .B(_19204_),
    .C(_19195_),
    .X(_03915_));
 sky130_fd_sc_hd__or2_1 _22088_ (.A(_19139_),
    .B(_19162_),
    .X(_19205_));
 sky130_fd_sc_hd__nand2_1 _22089_ (.A(_19205_),
    .B(_19138_),
    .Y(_19206_));
 sky130_fd_sc_hd__and3_1 _22090_ (.A(_19206_),
    .B(_19189_),
    .C(_19203_),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_1 _22091_ (.A(_19162_),
    .B(_19139_),
    .Y(_19207_));
 sky130_fd_sc_hd__and3_1 _22092_ (.A(_19205_),
    .B(_19189_),
    .C(_19207_),
    .X(_03913_));
 sky130_fd_sc_hd__nand2_1 _22093_ (.A(_19136_),
    .B(_19137_),
    .Y(_19208_));
 sky130_fd_sc_hd__nor2_1 _22094_ (.A(_19160_),
    .B(_19208_),
    .Y(_19209_));
 sky130_fd_sc_hd__nand2_1 _22095_ (.A(_19209_),
    .B(\count_instr[44] ),
    .Y(_19210_));
 sky130_fd_sc_hd__nor2_2 _22096_ (.A(_19142_),
    .B(_19210_),
    .Y(_19211_));
 sky130_fd_sc_hd__a21o_1 _22097_ (.A1(_19211_),
    .A2(\count_instr[46] ),
    .B1(\count_instr[47] ),
    .X(_19212_));
 sky130_fd_sc_hd__clkbuf_2 _22098_ (.A(_18542_),
    .X(_19213_));
 sky130_fd_sc_hd__and3_1 _22099_ (.A(_19212_),
    .B(_19213_),
    .C(_19162_),
    .X(_03912_));
 sky130_fd_sc_hd__o21ai_1 _22100_ (.A1(\count_instr[46] ),
    .A2(_19211_),
    .B1(_19175_),
    .Y(_19214_));
 sky130_fd_sc_hd__a21oi_1 _22101_ (.A1(\count_instr[46] ),
    .A2(_19211_),
    .B1(_19214_),
    .Y(_03911_));
 sky130_fd_sc_hd__or2_1 _22102_ (.A(_18793_),
    .B(_19211_),
    .X(_19215_));
 sky130_fd_sc_hd__a21oi_1 _22103_ (.A1(_19142_),
    .A2(_19210_),
    .B1(_19215_),
    .Y(_03910_));
 sky130_vsdinv _22104_ (.A(_19209_),
    .Y(_19216_));
 sky130_fd_sc_hd__nand2_1 _22105_ (.A(_19216_),
    .B(_19143_),
    .Y(_19217_));
 sky130_fd_sc_hd__and3_1 _22106_ (.A(_19217_),
    .B(_19213_),
    .C(_19210_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _22107_ (.A(_19208_),
    .B(_19160_),
    .Y(_19218_));
 sky130_fd_sc_hd__and3_1 _22108_ (.A(_19216_),
    .B(_19213_),
    .C(_19218_),
    .X(_03908_));
 sky130_fd_sc_hd__nor2_2 _22109_ (.A(_19093_),
    .B(_19135_),
    .Y(_19219_));
 sky130_fd_sc_hd__clkbuf_2 _22110_ (.A(\count_instr[37] ),
    .X(_19220_));
 sky130_fd_sc_hd__and3_1 _22111_ (.A(_19094_),
    .B(\count_instr[40] ),
    .C(_19220_),
    .X(_19221_));
 sky130_fd_sc_hd__a31o_1 _22112_ (.A1(_19219_),
    .A2(\count_instr[41] ),
    .A3(_19221_),
    .B1(\count_instr[42] ),
    .X(_19222_));
 sky130_fd_sc_hd__and3_1 _22113_ (.A(_19222_),
    .B(_19213_),
    .C(_19208_),
    .X(_03907_));
 sky130_vsdinv _22114_ (.A(\count_instr[41] ),
    .Y(_19223_));
 sky130_vsdinv _22115_ (.A(\count_instr[40] ),
    .Y(_19224_));
 sky130_vsdinv _22116_ (.A(_19136_),
    .Y(_19225_));
 sky130_fd_sc_hd__clkbuf_2 _22117_ (.A(_19219_),
    .X(_19226_));
 sky130_fd_sc_hd__a21o_1 _22118_ (.A1(_19226_),
    .A2(_19221_),
    .B1(\count_instr[41] ),
    .X(_19227_));
 sky130_fd_sc_hd__o311a_1 _22119_ (.A1(_19223_),
    .A2(_19224_),
    .A3(_19225_),
    .B1(_18543_),
    .C1(_19227_),
    .X(_03906_));
 sky130_fd_sc_hd__a221oi_2 _22120_ (.A1(_19226_),
    .A2(_19221_),
    .B1(_19225_),
    .B2(_19224_),
    .C1(_18794_),
    .Y(_03905_));
 sky130_fd_sc_hd__and3_1 _22121_ (.A(_19219_),
    .B(\count_instr[38] ),
    .C(_19220_),
    .X(_19228_));
 sky130_fd_sc_hd__or2_1 _22122_ (.A(\count_instr[39] ),
    .B(_19228_),
    .X(_19229_));
 sky130_fd_sc_hd__and3_1 _22123_ (.A(_19229_),
    .B(_19213_),
    .C(_19225_),
    .X(_03904_));
 sky130_fd_sc_hd__a21oi_1 _22124_ (.A1(_19226_),
    .A2(_19220_),
    .B1(\count_instr[38] ),
    .Y(_19230_));
 sky130_fd_sc_hd__nor3_1 _22125_ (.A(_19179_),
    .B(_19230_),
    .C(_19228_),
    .Y(_03903_));
 sky130_fd_sc_hd__o21ai_1 _22126_ (.A1(_19220_),
    .A2(_19226_),
    .B1(_19175_),
    .Y(_19231_));
 sky130_fd_sc_hd__a21oi_1 _22127_ (.A1(_19220_),
    .A2(_19226_),
    .B1(_19231_),
    .Y(_03902_));
 sky130_vsdinv _22128_ (.A(\count_instr[35] ),
    .Y(_19232_));
 sky130_vsdinv _22129_ (.A(\count_instr[34] ),
    .Y(_19233_));
 sky130_vsdinv _22130_ (.A(\count_instr[33] ),
    .Y(_19234_));
 sky130_fd_sc_hd__nand2_1 _22131_ (.A(_19126_),
    .B(\count_instr[27] ),
    .Y(_19235_));
 sky130_fd_sc_hd__nor2_1 _22132_ (.A(_19132_),
    .B(_19235_),
    .Y(_19236_));
 sky130_fd_sc_hd__nand2_1 _22133_ (.A(_19236_),
    .B(\count_instr[32] ),
    .Y(_19237_));
 sky130_fd_sc_hd__or2_1 _22134_ (.A(_19234_),
    .B(_19237_),
    .X(_19238_));
 sky130_fd_sc_hd__or3_1 _22135_ (.A(_19232_),
    .B(_19233_),
    .C(_19238_),
    .X(_19239_));
 sky130_vsdinv _22136_ (.A(\count_instr[36] ),
    .Y(_19240_));
 sky130_fd_sc_hd__or2_1 _22137_ (.A(_18793_),
    .B(_19226_),
    .X(_19241_));
 sky130_fd_sc_hd__a21oi_1 _22138_ (.A1(_19239_),
    .A2(_19240_),
    .B1(_19241_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _22139_ (.A(_19135_),
    .B(_19232_),
    .Y(_19242_));
 sky130_fd_sc_hd__and3_1 _22140_ (.A(_19239_),
    .B(_19213_),
    .C(_19242_),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_1 _22141_ (.A(_19238_),
    .B(_19233_),
    .Y(_19243_));
 sky130_fd_sc_hd__buf_2 _22142_ (.A(_18541_),
    .X(_19244_));
 sky130_fd_sc_hd__clkbuf_2 _22143_ (.A(_19244_),
    .X(_19245_));
 sky130_fd_sc_hd__and3_1 _22144_ (.A(_19243_),
    .B(_19245_),
    .C(_19135_),
    .X(_03899_));
 sky130_fd_sc_hd__nand2_1 _22145_ (.A(_19237_),
    .B(_19234_),
    .Y(_19246_));
 sky130_fd_sc_hd__and3_1 _22146_ (.A(_19238_),
    .B(_19245_),
    .C(_19246_),
    .X(_03898_));
 sky130_fd_sc_hd__or2_1 _22147_ (.A(\count_instr[32] ),
    .B(_19236_),
    .X(_19247_));
 sky130_fd_sc_hd__and3_1 _22148_ (.A(_19247_),
    .B(_19245_),
    .C(_19237_),
    .X(_03897_));
 sky130_fd_sc_hd__or2_2 _22149_ (.A(_19131_),
    .B(_19235_),
    .X(_19248_));
 sky130_fd_sc_hd__or3_1 _22150_ (.A(_19129_),
    .B(_19130_),
    .C(_19248_),
    .X(_19249_));
 sky130_fd_sc_hd__or2_1 _22151_ (.A(_18793_),
    .B(_19236_),
    .X(_19250_));
 sky130_fd_sc_hd__a21oi_1 _22152_ (.A1(_19249_),
    .A2(_19128_),
    .B1(_19250_),
    .Y(_03896_));
 sky130_fd_sc_hd__nor2_1 _22153_ (.A(_19130_),
    .B(_19248_),
    .Y(_19251_));
 sky130_fd_sc_hd__o211a_1 _22154_ (.A1(\count_instr[30] ),
    .A2(_19251_),
    .B1(_19090_),
    .C1(_19249_),
    .X(_03895_));
 sky130_fd_sc_hd__buf_2 _22155_ (.A(_18756_),
    .X(_19252_));
 sky130_fd_sc_hd__or2_1 _22156_ (.A(_19252_),
    .B(_19251_),
    .X(_19253_));
 sky130_fd_sc_hd__a21oi_1 _22157_ (.A1(_19130_),
    .A2(_19248_),
    .B1(_19253_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _22158_ (.A(_19235_),
    .B(_19131_),
    .Y(_19254_));
 sky130_fd_sc_hd__and3_1 _22159_ (.A(_19248_),
    .B(_19245_),
    .C(_19254_),
    .X(_03893_));
 sky130_fd_sc_hd__or2_1 _22160_ (.A(\count_instr[27] ),
    .B(_19126_),
    .X(_19255_));
 sky130_fd_sc_hd__and3_1 _22161_ (.A(_19255_),
    .B(_19245_),
    .C(_19235_),
    .X(_03892_));
 sky130_fd_sc_hd__nor2_1 _22162_ (.A(_19096_),
    .B(_19125_),
    .Y(_19256_));
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_18843_),
    .B(_19126_),
    .Y(_19257_));
 sky130_fd_sc_hd__o21a_1 _22164_ (.A1(\count_instr[26] ),
    .A2(_19256_),
    .B1(_19257_),
    .X(_03891_));
 sky130_fd_sc_hd__or2_1 _22165_ (.A(_19252_),
    .B(_19256_),
    .X(_19258_));
 sky130_fd_sc_hd__a21oi_1 _22166_ (.A1(_19096_),
    .A2(_19125_),
    .B1(_19258_),
    .Y(_03890_));
 sky130_vsdinv _22167_ (.A(\count_instr[23] ),
    .Y(_19259_));
 sky130_vsdinv _22168_ (.A(\count_instr[22] ),
    .Y(_19260_));
 sky130_fd_sc_hd__nand2_1 _22169_ (.A(_19120_),
    .B(\count_instr[19] ),
    .Y(_19261_));
 sky130_fd_sc_hd__nor2_1 _22170_ (.A(_19121_),
    .B(_19261_),
    .Y(_19262_));
 sky130_fd_sc_hd__nand2_1 _22171_ (.A(_19262_),
    .B(\count_instr[21] ),
    .Y(_19263_));
 sky130_fd_sc_hd__or3_1 _22172_ (.A(_19259_),
    .B(_19260_),
    .C(_19263_),
    .X(_19264_));
 sky130_vsdinv _22173_ (.A(\count_instr[24] ),
    .Y(_19265_));
 sky130_fd_sc_hd__nand2_1 _22174_ (.A(_19264_),
    .B(_19265_),
    .Y(_19266_));
 sky130_fd_sc_hd__and3_1 _22175_ (.A(_19266_),
    .B(_19245_),
    .C(_19125_),
    .X(_03889_));
 sky130_fd_sc_hd__nor2_1 _22176_ (.A(_19260_),
    .B(_19263_),
    .Y(_19267_));
 sky130_fd_sc_hd__o211a_1 _22177_ (.A1(\count_instr[23] ),
    .A2(_19267_),
    .B1(_19090_),
    .C1(_19264_),
    .X(_03888_));
 sky130_fd_sc_hd__or2_1 _22178_ (.A(_19252_),
    .B(_19267_),
    .X(_19268_));
 sky130_fd_sc_hd__a21oi_1 _22179_ (.A1(_19260_),
    .A2(_19263_),
    .B1(_19268_),
    .Y(_03887_));
 sky130_fd_sc_hd__or2_1 _22180_ (.A(\count_instr[21] ),
    .B(_19262_),
    .X(_19269_));
 sky130_fd_sc_hd__buf_2 _22181_ (.A(_19244_),
    .X(_19270_));
 sky130_fd_sc_hd__and3_1 _22182_ (.A(_19269_),
    .B(_19270_),
    .C(_19263_),
    .X(_03886_));
 sky130_fd_sc_hd__or2_1 _22183_ (.A(_19252_),
    .B(_19262_),
    .X(_19271_));
 sky130_fd_sc_hd__a21oi_1 _22184_ (.A1(_19121_),
    .A2(_19261_),
    .B1(_19271_),
    .Y(_03885_));
 sky130_fd_sc_hd__or2_1 _22185_ (.A(\count_instr[19] ),
    .B(_19120_),
    .X(_19272_));
 sky130_fd_sc_hd__and3_1 _22186_ (.A(_19272_),
    .B(_19270_),
    .C(_19261_),
    .X(_03884_));
 sky130_vsdinv _22187_ (.A(\count_instr[17] ),
    .Y(_19273_));
 sky130_vsdinv _22188_ (.A(_19119_),
    .Y(_19274_));
 sky130_fd_sc_hd__nor2_1 _22189_ (.A(_19273_),
    .B(_19274_),
    .Y(_19275_));
 sky130_fd_sc_hd__nor2_1 _22190_ (.A(_18843_),
    .B(_19120_),
    .Y(_19276_));
 sky130_fd_sc_hd__o21a_1 _22191_ (.A1(\count_instr[18] ),
    .A2(_19275_),
    .B1(_19276_),
    .X(_03883_));
 sky130_fd_sc_hd__o21ai_1 _22192_ (.A1(\count_instr[17] ),
    .A2(_19119_),
    .B1(_19175_),
    .Y(_19277_));
 sky130_fd_sc_hd__nor2_1 _22193_ (.A(_19277_),
    .B(_19275_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _22194_ (.A(_19118_),
    .B(_19097_),
    .Y(_19278_));
 sky130_fd_sc_hd__and3_1 _22195_ (.A(_19274_),
    .B(_19270_),
    .C(_19278_),
    .X(_03881_));
 sky130_fd_sc_hd__or2_1 _22196_ (.A(\count_instr[15] ),
    .B(_19117_),
    .X(_19279_));
 sky130_fd_sc_hd__and3_1 _22197_ (.A(_19279_),
    .B(_19270_),
    .C(_19118_),
    .X(_03880_));
 sky130_fd_sc_hd__or2_1 _22198_ (.A(_19252_),
    .B(_19117_),
    .X(_19280_));
 sky130_fd_sc_hd__a21oi_1 _22199_ (.A1(_19098_),
    .A2(_19116_),
    .B1(_19280_),
    .Y(_03879_));
 sky130_fd_sc_hd__nor2_2 _22200_ (.A(_19115_),
    .B(_18663_),
    .Y(_19281_));
 sky130_fd_sc_hd__o211a_1 _22201_ (.A1(\count_instr[13] ),
    .A2(_19281_),
    .B1(_19090_),
    .C1(_19116_),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_1 _22202_ (.A(_18664_),
    .B(\count_instr[0] ),
    .Y(_19282_));
 sky130_fd_sc_hd__or2_1 _22203_ (.A(_19110_),
    .B(_19282_),
    .X(_19283_));
 sky130_fd_sc_hd__or2_1 _22204_ (.A(_19109_),
    .B(_19283_),
    .X(_19284_));
 sky130_fd_sc_hd__or2_1 _22205_ (.A(_19099_),
    .B(_19284_),
    .X(_19285_));
 sky130_fd_sc_hd__nor2_1 _22206_ (.A(_19108_),
    .B(_19285_),
    .Y(_19286_));
 sky130_fd_sc_hd__nand2_1 _22207_ (.A(_19286_),
    .B(\count_instr[6] ),
    .Y(_19287_));
 sky130_fd_sc_hd__nor2_1 _22208_ (.A(_19102_),
    .B(_19287_),
    .Y(_19288_));
 sky130_fd_sc_hd__nand2_1 _22209_ (.A(_19288_),
    .B(\count_instr[8] ),
    .Y(_19289_));
 sky130_fd_sc_hd__nor2_1 _22210_ (.A(_19106_),
    .B(_19289_),
    .Y(_19290_));
 sky130_fd_sc_hd__nand2_1 _22211_ (.A(_19290_),
    .B(\count_instr[10] ),
    .Y(_19291_));
 sky130_fd_sc_hd__or2_1 _22212_ (.A(_19101_),
    .B(_19291_),
    .X(_19292_));
 sky130_fd_sc_hd__a211oi_2 _22213_ (.A1(_19292_),
    .A2(_19100_),
    .B1(_18794_),
    .C1(_19281_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _22214_ (.A(_19291_),
    .B(_19101_),
    .Y(_19293_));
 sky130_fd_sc_hd__and3_1 _22215_ (.A(_19292_),
    .B(_19270_),
    .C(_19293_),
    .X(_03876_));
 sky130_vsdinv _22216_ (.A(_19290_),
    .Y(_19294_));
 sky130_fd_sc_hd__nand2_1 _22217_ (.A(_19294_),
    .B(_19105_),
    .Y(_19295_));
 sky130_fd_sc_hd__and3_1 _22218_ (.A(_19295_),
    .B(_19270_),
    .C(_19291_),
    .X(_03875_));
 sky130_fd_sc_hd__buf_1 _22219_ (.A(_19244_),
    .X(_19296_));
 sky130_fd_sc_hd__nand2_1 _22220_ (.A(_19289_),
    .B(_19106_),
    .Y(_19297_));
 sky130_fd_sc_hd__and3_1 _22221_ (.A(_19294_),
    .B(_19296_),
    .C(_19297_),
    .X(_03874_));
 sky130_vsdinv _22222_ (.A(_19288_),
    .Y(_19298_));
 sky130_fd_sc_hd__nand2_1 _22223_ (.A(_19298_),
    .B(_19107_),
    .Y(_19299_));
 sky130_fd_sc_hd__and3_1 _22224_ (.A(_19299_),
    .B(_19296_),
    .C(_19289_),
    .X(_03873_));
 sky130_fd_sc_hd__nand2_1 _22225_ (.A(_19287_),
    .B(_19102_),
    .Y(_19300_));
 sky130_fd_sc_hd__and3_1 _22226_ (.A(_19298_),
    .B(_19296_),
    .C(_19300_),
    .X(_03872_));
 sky130_vsdinv _22227_ (.A(_19286_),
    .Y(_19301_));
 sky130_fd_sc_hd__nand2_1 _22228_ (.A(_19301_),
    .B(_19103_),
    .Y(_19302_));
 sky130_fd_sc_hd__and3_1 _22229_ (.A(_19302_),
    .B(_19296_),
    .C(_19287_),
    .X(_03871_));
 sky130_fd_sc_hd__nand2_1 _22230_ (.A(_19285_),
    .B(_19108_),
    .Y(_19303_));
 sky130_fd_sc_hd__and3_1 _22231_ (.A(_19301_),
    .B(_19296_),
    .C(_19303_),
    .X(_03870_));
 sky130_vsdinv _22232_ (.A(\count_instr[3] ),
    .Y(_19304_));
 sky130_fd_sc_hd__or2_1 _22233_ (.A(_19304_),
    .B(_19284_),
    .X(_19305_));
 sky130_vsdinv _22234_ (.A(\count_instr[4] ),
    .Y(_19306_));
 sky130_fd_sc_hd__nand2_1 _22235_ (.A(_19305_),
    .B(_19306_),
    .Y(_19307_));
 sky130_fd_sc_hd__and3_1 _22236_ (.A(_19307_),
    .B(_19296_),
    .C(_19285_),
    .X(_03869_));
 sky130_fd_sc_hd__buf_2 _22237_ (.A(_19244_),
    .X(_19308_));
 sky130_fd_sc_hd__nand2_1 _22238_ (.A(_19284_),
    .B(_19304_),
    .Y(_19309_));
 sky130_fd_sc_hd__and3_1 _22239_ (.A(_19305_),
    .B(_19308_),
    .C(_19309_),
    .X(_03868_));
 sky130_fd_sc_hd__nand2_1 _22240_ (.A(_19283_),
    .B(_19109_),
    .Y(_19310_));
 sky130_fd_sc_hd__and3_1 _22241_ (.A(_19284_),
    .B(_19308_),
    .C(_19310_),
    .X(_03867_));
 sky130_fd_sc_hd__nand2_1 _22242_ (.A(_19282_),
    .B(_19110_),
    .Y(_19311_));
 sky130_fd_sc_hd__and3_1 _22243_ (.A(_19283_),
    .B(_19308_),
    .C(_19311_),
    .X(_03866_));
 sky130_fd_sc_hd__nand2_1 _22244_ (.A(_18663_),
    .B(_19111_),
    .Y(_19312_));
 sky130_fd_sc_hd__and3_1 _22245_ (.A(_19282_),
    .B(_19308_),
    .C(_19312_),
    .X(_03865_));
 sky130_fd_sc_hd__and3_1 _22246_ (.A(_18750_),
    .B(_18552_),
    .C(_18775_),
    .X(_19313_));
 sky130_fd_sc_hd__buf_2 _22247_ (.A(_19313_),
    .X(_19314_));
 sky130_fd_sc_hd__clkbuf_2 _22248_ (.A(_19314_),
    .X(_19315_));
 sky130_fd_sc_hd__clkbuf_2 _22249_ (.A(_18706_),
    .X(_19316_));
 sky130_fd_sc_hd__clkbuf_4 _22250_ (.A(_19316_),
    .X(_19317_));
 sky130_vsdinv _22251_ (.A(_19313_),
    .Y(_19318_));
 sky130_fd_sc_hd__clkbuf_2 _22252_ (.A(_19318_),
    .X(_19319_));
 sky130_fd_sc_hd__clkbuf_2 _22253_ (.A(_19319_),
    .X(_19320_));
 sky130_fd_sc_hd__a21o_1 _22254_ (.A1(_19317_),
    .A2(_18641_),
    .B1(_19320_),
    .X(_19321_));
 sky130_fd_sc_hd__o211a_1 _22255_ (.A1(net126),
    .A2(_19315_),
    .B1(_19090_),
    .C1(_19321_),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_2 _22256_ (.A(_19048_),
    .X(_19322_));
 sky130_fd_sc_hd__a21o_1 _22257_ (.A1(_19317_),
    .A2(_18643_),
    .B1(_19320_),
    .X(_19323_));
 sky130_fd_sc_hd__o211a_1 _22258_ (.A1(net125),
    .A2(_19315_),
    .B1(_19322_),
    .C1(_19323_),
    .X(_03863_));
 sky130_fd_sc_hd__buf_2 _22259_ (.A(_18707_),
    .X(_19324_));
 sky130_fd_sc_hd__buf_2 _22260_ (.A(_19318_),
    .X(_19325_));
 sky130_fd_sc_hd__a31o_1 _22261_ (.A1(_18637_),
    .A2(_19324_),
    .A3(\irq_pending[29] ),
    .B1(_19325_),
    .X(_19326_));
 sky130_fd_sc_hd__o211a_1 _22262_ (.A1(net123),
    .A2(_19315_),
    .B1(_19322_),
    .C1(_19326_),
    .X(_03862_));
 sky130_fd_sc_hd__a21o_1 _22263_ (.A1(_19317_),
    .A2(_18639_),
    .B1(_19320_),
    .X(_19327_));
 sky130_fd_sc_hd__o211a_1 _22264_ (.A1(net122),
    .A2(_19315_),
    .B1(_19322_),
    .C1(_19327_),
    .X(_03861_));
 sky130_fd_sc_hd__a21o_1 _22265_ (.A1(_19317_),
    .A2(_18611_),
    .B1(_19320_),
    .X(_19328_));
 sky130_fd_sc_hd__o211a_1 _22266_ (.A1(net121),
    .A2(_19315_),
    .B1(_19322_),
    .C1(_19328_),
    .X(_03860_));
 sky130_fd_sc_hd__a21o_1 _22267_ (.A1(_19317_),
    .A2(_18612_),
    .B1(_19320_),
    .X(_19329_));
 sky130_fd_sc_hd__o211a_1 _22268_ (.A1(net120),
    .A2(_19315_),
    .B1(_19322_),
    .C1(_19329_),
    .X(_03859_));
 sky130_fd_sc_hd__clkbuf_2 _22269_ (.A(_19314_),
    .X(_19330_));
 sky130_fd_sc_hd__a31o_1 _22270_ (.A1(_18613_),
    .A2(_19324_),
    .A3(\irq_pending[25] ),
    .B1(_19325_),
    .X(_19331_));
 sky130_fd_sc_hd__o211a_1 _22271_ (.A1(net119),
    .A2(_19330_),
    .B1(_19322_),
    .C1(_19331_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_2 _22272_ (.A(_19048_),
    .X(_19332_));
 sky130_fd_sc_hd__buf_2 _22273_ (.A(_18707_),
    .X(_19333_));
 sky130_fd_sc_hd__a31o_1 _22274_ (.A1(_18614_),
    .A2(_19333_),
    .A3(\irq_pending[24] ),
    .B1(_19325_),
    .X(_19334_));
 sky130_fd_sc_hd__o211a_1 _22275_ (.A1(net118),
    .A2(_19330_),
    .B1(_19332_),
    .C1(_19334_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_2 _22276_ (.A(_18706_),
    .X(_19335_));
 sky130_fd_sc_hd__buf_2 _22277_ (.A(_19335_),
    .X(_19336_));
 sky130_fd_sc_hd__a21o_1 _22278_ (.A1(_19336_),
    .A2(_18618_),
    .B1(_19320_),
    .X(_19337_));
 sky130_fd_sc_hd__o211a_1 _22279_ (.A1(net117),
    .A2(_19330_),
    .B1(_19332_),
    .C1(_19337_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_2 _22280_ (.A(_19319_),
    .X(_19338_));
 sky130_fd_sc_hd__a21o_1 _22281_ (.A1(_19336_),
    .A2(_18619_),
    .B1(_19338_),
    .X(_19339_));
 sky130_fd_sc_hd__o211a_1 _22282_ (.A1(net116),
    .A2(_19330_),
    .B1(_19332_),
    .C1(_19339_),
    .X(_03855_));
 sky130_fd_sc_hd__a31o_1 _22283_ (.A1(_18620_),
    .A2(_19333_),
    .A3(\irq_pending[21] ),
    .B1(_19325_),
    .X(_19340_));
 sky130_fd_sc_hd__o211a_1 _22284_ (.A1(net115),
    .A2(_19330_),
    .B1(_19332_),
    .C1(_19340_),
    .X(_03854_));
 sky130_fd_sc_hd__buf_2 _22285_ (.A(_19319_),
    .X(_19341_));
 sky130_fd_sc_hd__a31o_1 _22286_ (.A1(_18621_),
    .A2(_19333_),
    .A3(\irq_pending[20] ),
    .B1(_19341_),
    .X(_19342_));
 sky130_fd_sc_hd__o211a_1 _22287_ (.A1(net114),
    .A2(_19330_),
    .B1(_19332_),
    .C1(_19342_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_2 _22288_ (.A(_19314_),
    .X(_19343_));
 sky130_fd_sc_hd__a21o_1 _22289_ (.A1(_19336_),
    .A2(_18607_),
    .B1(_19338_),
    .X(_19344_));
 sky130_fd_sc_hd__o211a_1 _22290_ (.A1(net112),
    .A2(_19343_),
    .B1(_19332_),
    .C1(_19344_),
    .X(_03852_));
 sky130_fd_sc_hd__buf_2 _22291_ (.A(_18542_),
    .X(_19345_));
 sky130_fd_sc_hd__a21o_1 _22292_ (.A1(_19336_),
    .A2(_18609_),
    .B1(_19338_),
    .X(_19346_));
 sky130_fd_sc_hd__o211a_1 _22293_ (.A1(net111),
    .A2(_19343_),
    .B1(_19345_),
    .C1(_19346_),
    .X(_03851_));
 sky130_fd_sc_hd__a31o_1 _22294_ (.A1(_18603_),
    .A2(_19333_),
    .A3(\irq_pending[17] ),
    .B1(_19341_),
    .X(_19347_));
 sky130_fd_sc_hd__o211a_1 _22295_ (.A1(net110),
    .A2(_19343_),
    .B1(_19345_),
    .C1(_19347_),
    .X(_03850_));
 sky130_fd_sc_hd__a21o_1 _22296_ (.A1(_19336_),
    .A2(_18605_),
    .B1(_19338_),
    .X(_19348_));
 sky130_fd_sc_hd__o211a_1 _22297_ (.A1(net109),
    .A2(_19343_),
    .B1(_19345_),
    .C1(_19348_),
    .X(_03849_));
 sky130_fd_sc_hd__a21o_1 _22298_ (.A1(_19336_),
    .A2(_18649_),
    .B1(_19338_),
    .X(_19349_));
 sky130_fd_sc_hd__o211a_1 _22299_ (.A1(net108),
    .A2(_19343_),
    .B1(_19345_),
    .C1(_19349_),
    .X(_03848_));
 sky130_fd_sc_hd__clkbuf_2 _22300_ (.A(_19335_),
    .X(_19350_));
 sky130_fd_sc_hd__a21o_1 _22301_ (.A1(_19350_),
    .A2(_18651_),
    .B1(_19338_),
    .X(_19351_));
 sky130_fd_sc_hd__o211a_1 _22302_ (.A1(net107),
    .A2(_19343_),
    .B1(_19345_),
    .C1(_19351_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_2 _22303_ (.A(_19314_),
    .X(_19352_));
 sky130_fd_sc_hd__a31o_1 _22304_ (.A1(_18645_),
    .A2(_19333_),
    .A3(\irq_pending[13] ),
    .B1(_19341_),
    .X(_19353_));
 sky130_fd_sc_hd__o211a_1 _22305_ (.A1(net106),
    .A2(_19352_),
    .B1(_19345_),
    .C1(_19353_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_2 _22306_ (.A(_18542_),
    .X(_19354_));
 sky130_fd_sc_hd__clkbuf_2 _22307_ (.A(_19319_),
    .X(_19355_));
 sky130_fd_sc_hd__a21o_1 _22308_ (.A1(_19350_),
    .A2(_18647_),
    .B1(_19355_),
    .X(_19356_));
 sky130_fd_sc_hd__o211a_1 _22309_ (.A1(net105),
    .A2(_19352_),
    .B1(_19354_),
    .C1(_19356_),
    .X(_03845_));
 sky130_fd_sc_hd__a21o_1 _22310_ (.A1(_19350_),
    .A2(_18625_),
    .B1(_19355_),
    .X(_19357_));
 sky130_fd_sc_hd__o211a_1 _22311_ (.A1(net104),
    .A2(_19352_),
    .B1(_19354_),
    .C1(_19357_),
    .X(_03844_));
 sky130_fd_sc_hd__a21o_1 _22312_ (.A1(_19350_),
    .A2(_18626_),
    .B1(_19355_),
    .X(_19358_));
 sky130_fd_sc_hd__o211a_1 _22313_ (.A1(net103),
    .A2(_19352_),
    .B1(_19354_),
    .C1(_19358_),
    .X(_03843_));
 sky130_fd_sc_hd__a31o_1 _22314_ (.A1(_18627_),
    .A2(_19333_),
    .A3(\irq_pending[9] ),
    .B1(_19341_),
    .X(_19359_));
 sky130_fd_sc_hd__o211a_1 _22315_ (.A1(net133),
    .A2(_19352_),
    .B1(_19354_),
    .C1(_19359_),
    .X(_03842_));
 sky130_fd_sc_hd__buf_2 _22316_ (.A(_18707_),
    .X(_19360_));
 sky130_fd_sc_hd__a31o_1 _22317_ (.A1(_18628_),
    .A2(_19360_),
    .A3(\irq_pending[8] ),
    .B1(_19341_),
    .X(_19361_));
 sky130_fd_sc_hd__o211a_1 _22318_ (.A1(net132),
    .A2(_19352_),
    .B1(_19354_),
    .C1(_19361_),
    .X(_03841_));
 sky130_fd_sc_hd__clkbuf_2 _22319_ (.A(_19313_),
    .X(_19362_));
 sky130_fd_sc_hd__a21o_1 _22320_ (.A1(_19350_),
    .A2(_18631_),
    .B1(_19355_),
    .X(_19363_));
 sky130_fd_sc_hd__o211a_1 _22321_ (.A1(net131),
    .A2(_19362_),
    .B1(_19354_),
    .C1(_19363_),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_2 _22322_ (.A(_18542_),
    .X(_19364_));
 sky130_fd_sc_hd__a21o_1 _22323_ (.A1(_19350_),
    .A2(_18632_),
    .B1(_19355_),
    .X(_19365_));
 sky130_fd_sc_hd__o211a_1 _22324_ (.A1(net130),
    .A2(_19362_),
    .B1(_19364_),
    .C1(_19365_),
    .X(_03839_));
 sky130_fd_sc_hd__a31o_1 _22325_ (.A1(_18633_),
    .A2(_19360_),
    .A3(\irq_pending[5] ),
    .B1(_19341_),
    .X(_19366_));
 sky130_fd_sc_hd__o211a_1 _22326_ (.A1(net129),
    .A2(_19362_),
    .B1(_19364_),
    .C1(_19366_),
    .X(_03838_));
 sky130_fd_sc_hd__a31o_1 _22327_ (.A1(_18634_),
    .A2(_19360_),
    .A3(\irq_pending[4] ),
    .B1(_19319_),
    .X(_19367_));
 sky130_fd_sc_hd__o211a_1 _22328_ (.A1(net128),
    .A2(_19362_),
    .B1(_19364_),
    .C1(_19367_),
    .X(_03837_));
 sky130_fd_sc_hd__a21o_1 _22329_ (.A1(_19324_),
    .A2(_18601_),
    .B1(_19355_),
    .X(_19368_));
 sky130_fd_sc_hd__o211a_1 _22330_ (.A1(net127),
    .A2(_19362_),
    .B1(_19364_),
    .C1(_19368_),
    .X(_03836_));
 sky130_fd_sc_hd__a31o_1 _22331_ (.A1(_18595_),
    .A2(_19360_),
    .A3(\irq_pending[2] ),
    .B1(_19319_),
    .X(_19369_));
 sky130_fd_sc_hd__o211a_1 _22332_ (.A1(net124),
    .A2(_19362_),
    .B1(_19364_),
    .C1(_19369_),
    .X(_03835_));
 sky130_fd_sc_hd__a21o_1 _22333_ (.A1(_19324_),
    .A2(_18599_),
    .B1(_19325_),
    .X(_19370_));
 sky130_fd_sc_hd__o211a_1 _22334_ (.A1(net113),
    .A2(_19314_),
    .B1(_19364_),
    .C1(_19370_),
    .X(_03834_));
 sky130_fd_sc_hd__a21o_1 _22335_ (.A1(_19324_),
    .A2(_18597_),
    .B1(_19325_),
    .X(_19371_));
 sky130_fd_sc_hd__o211a_1 _22336_ (.A1(net102),
    .A2(_19314_),
    .B1(_19195_),
    .C1(_19371_),
    .X(_03833_));
 sky130_fd_sc_hd__nor2_4 _22337_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_vsdinv _22338_ (.A(_00311_),
    .Y(_19372_));
 sky130_fd_sc_hd__nor2_2 _22339_ (.A(_18743_),
    .B(_18764_),
    .Y(_19373_));
 sky130_vsdinv _22340_ (.A(_19373_),
    .Y(_19374_));
 sky130_fd_sc_hd__or3_4 _22341_ (.A(\pcpi_mul.active[1] ),
    .B(_19372_),
    .C(_19374_),
    .X(_19375_));
 sky130_fd_sc_hd__nand2_1 _22342_ (.A(_19374_),
    .B(net370),
    .Y(_19376_));
 sky130_fd_sc_hd__a21oi_1 _22343_ (.A1(_19375_),
    .A2(_19376_),
    .B1(_19179_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _22344_ (.A(_18564_),
    .B(_00290_),
    .Y(_19377_));
 sky130_fd_sc_hd__a21bo_1 _22345_ (.A1(_18560_),
    .A2(_18528_),
    .B1_N(net237),
    .X(_19378_));
 sky130_fd_sc_hd__a21o_1 _22346_ (.A1(_19377_),
    .A2(_19378_),
    .B1(net408),
    .X(_19379_));
 sky130_fd_sc_hd__or2b_1 _22347_ (.A(net521),
    .B_N(net237),
    .X(_19380_));
 sky130_fd_sc_hd__a21oi_1 _22348_ (.A1(_19379_),
    .A2(_19380_),
    .B1(_19179_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_4 _22349_ (.A(\irq_pending[25] ),
    .B(\irq_pending[24] ),
    .C(\irq_pending[27] ),
    .D(\irq_pending[26] ),
    .X(_19381_));
 sky130_fd_sc_hd__or4_4 _22350_ (.A(\irq_pending[21] ),
    .B(\irq_pending[20] ),
    .C(\irq_pending[23] ),
    .D(\irq_pending[22] ),
    .X(_19382_));
 sky130_fd_sc_hd__or4_4 _22351_ (.A(\irq_pending[17] ),
    .B(\irq_pending[16] ),
    .C(\irq_pending[19] ),
    .D(\irq_pending[18] ),
    .X(_19383_));
 sky130_fd_sc_hd__or4_4 _22352_ (.A(\irq_pending[29] ),
    .B(\irq_pending[28] ),
    .C(\irq_pending[31] ),
    .D(\irq_pending[30] ),
    .X(_19384_));
 sky130_fd_sc_hd__or4_4 _22353_ (.A(_19381_),
    .B(_19382_),
    .C(_19383_),
    .D(_19384_),
    .X(_19385_));
 sky130_fd_sc_hd__or4_4 _22354_ (.A(\irq_pending[9] ),
    .B(\irq_pending[8] ),
    .C(\irq_pending[11] ),
    .D(\irq_pending[10] ),
    .X(_19386_));
 sky130_fd_sc_hd__or4_4 _22355_ (.A(\irq_pending[5] ),
    .B(\irq_pending[4] ),
    .C(\irq_pending[7] ),
    .D(\irq_pending[6] ),
    .X(_19387_));
 sky130_fd_sc_hd__or4_4 _22356_ (.A(\irq_pending[1] ),
    .B(\irq_pending[0] ),
    .C(\irq_pending[3] ),
    .D(\irq_pending[2] ),
    .X(_19388_));
 sky130_fd_sc_hd__or4_4 _22357_ (.A(\irq_pending[13] ),
    .B(\irq_pending[12] ),
    .C(\irq_pending[15] ),
    .D(\irq_pending[14] ),
    .X(_19389_));
 sky130_fd_sc_hd__or4_4 _22358_ (.A(_19386_),
    .B(_19387_),
    .C(_19388_),
    .D(_19389_),
    .X(_19390_));
 sky130_fd_sc_hd__nor2_8 _22359_ (.A(_19385_),
    .B(_19390_),
    .Y(_02410_));
 sky130_fd_sc_hd__buf_6 _22360_ (.A(_18657_),
    .X(_00308_));
 sky130_fd_sc_hd__nor2_1 _22361_ (.A(_18532_),
    .B(_00308_),
    .Y(_19391_));
 sky130_fd_sc_hd__nand2_1 _22362_ (.A(_19391_),
    .B(_00309_),
    .Y(_19392_));
 sky130_vsdinv _22363_ (.A(_19392_),
    .Y(_19393_));
 sky130_fd_sc_hd__and3_1 _22364_ (.A(_19393_),
    .B(_19016_),
    .C(_02410_),
    .X(_03830_));
 sky130_fd_sc_hd__or4_4 _22365_ (.A(_18699_),
    .B(instr_sltu),
    .C(instr_slt),
    .D(_18726_),
    .X(_19394_));
 sky130_fd_sc_hd__buf_2 _22366_ (.A(_18904_),
    .X(_19395_));
 sky130_fd_sc_hd__and3_2 _22367_ (.A(_19394_),
    .B(_19308_),
    .C(_19395_),
    .X(_03829_));
 sky130_fd_sc_hd__and4_1 _22368_ (.A(_18772_),
    .B(_18540_),
    .C(_18964_),
    .D(_18777_),
    .X(_19396_));
 sky130_fd_sc_hd__buf_1 _22369_ (.A(_19396_),
    .X(_03828_));
 sky130_fd_sc_hd__nor2_1 _22370_ (.A(_18944_),
    .B(_18957_),
    .Y(_03827_));
 sky130_fd_sc_hd__clkbuf_4 _22371_ (.A(_18548_),
    .X(_19397_));
 sky130_fd_sc_hd__and2_1 _22372_ (.A(_19397_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_1 _22373_ (.A(_19397_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_1 _22374_ (.A(_19397_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_1 _22375_ (.A(_19397_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_1 _22376_ (.A(_19397_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_2 _22377_ (.A(_19175_),
    .X(_19398_));
 sky130_fd_sc_hd__and2_1 _22378_ (.A(_19398_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_1 _22379_ (.A(_19398_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__and2_1 _22380_ (.A(_19398_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _22381_ (.A(_19398_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__and2_1 _22382_ (.A(_19398_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_1 _22383_ (.A(_19398_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__buf_2 _22384_ (.A(_18547_),
    .X(_19399_));
 sky130_fd_sc_hd__clkbuf_2 _22385_ (.A(_19399_),
    .X(_19400_));
 sky130_fd_sc_hd__and2_1 _22386_ (.A(_19400_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _22387_ (.A(_19400_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__and2_1 _22388_ (.A(_19400_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_1 _22389_ (.A(_19400_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__and2_1 _22390_ (.A(_19400_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_1 _22391_ (.A(_19400_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_2 _22392_ (.A(_19399_),
    .X(_19401_));
 sky130_fd_sc_hd__and2_1 _22393_ (.A(_19401_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_1 _22394_ (.A(_19401_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_1 _22395_ (.A(_19401_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_1 _22396_ (.A(_19401_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_1 _22397_ (.A(_19401_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_1 _22398_ (.A(_19401_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_2 _22399_ (.A(_19399_),
    .X(_19402_));
 sky130_fd_sc_hd__and2_1 _22400_ (.A(_19402_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_1 _22401_ (.A(_19402_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_1 _22402_ (.A(_19402_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_1 _22403_ (.A(_19402_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__and2_1 _22404_ (.A(_19402_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_1 _22405_ (.A(_19402_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__clkbuf_2 _22406_ (.A(_19399_),
    .X(_19403_));
 sky130_fd_sc_hd__and2_1 _22407_ (.A(_19403_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_1 _22408_ (.A(_19403_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _22409_ (.A(_19403_),
    .B(_02411_),
    .X(_03795_));
 sky130_vsdinv _22410_ (.A(\count_cycle[56] ),
    .Y(_19404_));
 sky130_fd_sc_hd__nand2_1 _22411_ (.A(\count_cycle[54] ),
    .B(\count_cycle[55] ),
    .Y(_19405_));
 sky130_vsdinv _22412_ (.A(\count_cycle[51] ),
    .Y(_19406_));
 sky130_vsdinv _22413_ (.A(\count_cycle[52] ),
    .Y(_19407_));
 sky130_vsdinv _22414_ (.A(\count_cycle[53] ),
    .Y(_19408_));
 sky130_fd_sc_hd__or4_4 _22415_ (.A(_19405_),
    .B(_19406_),
    .C(_19407_),
    .D(_19408_),
    .X(_19409_));
 sky130_vsdinv _22416_ (.A(\count_cycle[38] ),
    .Y(_19410_));
 sky130_vsdinv _22417_ (.A(\count_cycle[39] ),
    .Y(_19411_));
 sky130_fd_sc_hd__nor2_1 _22418_ (.A(_19410_),
    .B(_19411_),
    .Y(_19412_));
 sky130_vsdinv _22419_ (.A(_19412_),
    .Y(_19413_));
 sky130_vsdinv _22420_ (.A(\count_cycle[40] ),
    .Y(_19414_));
 sky130_vsdinv _22421_ (.A(\count_cycle[41] ),
    .Y(_19415_));
 sky130_vsdinv _22422_ (.A(\count_cycle[42] ),
    .Y(_19416_));
 sky130_vsdinv _22423_ (.A(\count_cycle[43] ),
    .Y(_19417_));
 sky130_fd_sc_hd__or4_4 _22424_ (.A(_19414_),
    .B(_19415_),
    .C(_19416_),
    .D(_19417_),
    .X(_19418_));
 sky130_vsdinv _22425_ (.A(\count_cycle[33] ),
    .Y(_19419_));
 sky130_fd_sc_hd__inv_2 _22426_ (.A(\count_cycle[28] ),
    .Y(_02028_));
 sky130_fd_sc_hd__inv_2 _22427_ (.A(\count_cycle[29] ),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _22428_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_fd_sc_hd__inv_2 _22429_ (.A(\count_cycle[31] ),
    .Y(_02055_));
 sky130_fd_sc_hd__or4_4 _22430_ (.A(_02028_),
    .B(_02037_),
    .C(_02046_),
    .D(_02055_),
    .X(_19420_));
 sky130_fd_sc_hd__nor2_1 _22431_ (.A(_19419_),
    .B(_19420_),
    .Y(_19421_));
 sky130_vsdinv _22432_ (.A(_19421_),
    .Y(_19422_));
 sky130_fd_sc_hd__inv_2 _22433_ (.A(\count_cycle[22] ),
    .Y(_01974_));
 sky130_fd_sc_hd__inv_2 _22434_ (.A(\count_cycle[20] ),
    .Y(_01956_));
 sky130_fd_sc_hd__inv_2 _22435_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_fd_sc_hd__inv_2 _22436_ (.A(\count_cycle[16] ),
    .Y(_01920_));
 sky130_fd_sc_hd__inv_2 _22437_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__inv_2 _22438_ (.A(\count_cycle[13] ),
    .Y(_01885_));
 sky130_fd_sc_hd__inv_2 _22439_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_fd_sc_hd__inv_2 _22440_ (.A(\count_cycle[10] ),
    .Y(_01846_));
 sky130_fd_sc_hd__inv_2 _22441_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _22442_ (.A(\count_cycle[7] ),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _22443_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _22444_ (.A(\count_cycle[5] ),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_2 _22445_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_1 _22446_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .Y(_19423_));
 sky130_fd_sc_hd__inv_2 _22447_ (.A(\count_cycle[2] ),
    .Y(_01741_));
 sky130_fd_sc_hd__or2_1 _22448_ (.A(_19423_),
    .B(_01741_),
    .X(_19424_));
 sky130_fd_sc_hd__nor2_1 _22449_ (.A(_01754_),
    .B(_19424_),
    .Y(_19425_));
 sky130_fd_sc_hd__nand2_1 _22450_ (.A(_19425_),
    .B(\count_cycle[4] ),
    .Y(_19426_));
 sky130_fd_sc_hd__nor2_1 _22451_ (.A(_01780_),
    .B(_19426_),
    .Y(_19427_));
 sky130_fd_sc_hd__nand2_1 _22452_ (.A(_19427_),
    .B(\count_cycle[6] ),
    .Y(_19428_));
 sky130_fd_sc_hd__or3_1 _22453_ (.A(_01806_),
    .B(_01820_),
    .C(_19428_),
    .X(_19429_));
 sky130_fd_sc_hd__or2_1 _22454_ (.A(_01833_),
    .B(_19429_),
    .X(_19430_));
 sky130_fd_sc_hd__nor2_1 _22455_ (.A(_01846_),
    .B(_19430_),
    .Y(_19431_));
 sky130_fd_sc_hd__nand2_1 _22456_ (.A(_19431_),
    .B(\count_cycle[11] ),
    .Y(_19432_));
 sky130_fd_sc_hd__or2_1 _22457_ (.A(_01872_),
    .B(_19432_),
    .X(_19433_));
 sky130_fd_sc_hd__nor2_1 _22458_ (.A(_01885_),
    .B(_19433_),
    .Y(_19434_));
 sky130_fd_sc_hd__nand2_1 _22459_ (.A(_19434_),
    .B(\count_cycle[14] ),
    .Y(_19435_));
 sky130_fd_sc_hd__or2_1 _22460_ (.A(_01911_),
    .B(_19435_),
    .X(_19436_));
 sky130_fd_sc_hd__nor2_1 _22461_ (.A(_01920_),
    .B(_19436_),
    .Y(_19437_));
 sky130_fd_sc_hd__nand2_1 _22462_ (.A(_19437_),
    .B(\count_cycle[17] ),
    .Y(_19438_));
 sky130_fd_sc_hd__nor2_2 _22463_ (.A(_01938_),
    .B(_19438_),
    .Y(_19439_));
 sky130_fd_sc_hd__nand2_2 _22464_ (.A(_19439_),
    .B(\count_cycle[19] ),
    .Y(_19440_));
 sky130_fd_sc_hd__nor2_1 _22465_ (.A(_01956_),
    .B(_19440_),
    .Y(_19441_));
 sky130_fd_sc_hd__nand2_1 _22466_ (.A(_19441_),
    .B(\count_cycle[21] ),
    .Y(_19442_));
 sky130_fd_sc_hd__nor2_2 _22467_ (.A(_01974_),
    .B(_19442_),
    .Y(_19443_));
 sky130_fd_sc_hd__inv_2 _22468_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__inv_2 _22469_ (.A(\count_cycle[24] ),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _22470_ (.A(_01983_),
    .B(_01992_),
    .Y(_19444_));
 sky130_fd_sc_hd__and3_2 _22471_ (.A(_19443_),
    .B(\count_cycle[25] ),
    .C(_19444_),
    .X(_19445_));
 sky130_fd_sc_hd__inv_2 _22472_ (.A(\count_cycle[26] ),
    .Y(_02010_));
 sky130_fd_sc_hd__inv_2 _22473_ (.A(\count_cycle[27] ),
    .Y(_02019_));
 sky130_fd_sc_hd__nor2_2 _22474_ (.A(_02010_),
    .B(_02019_),
    .Y(_19446_));
 sky130_fd_sc_hd__nand3_4 _22475_ (.A(_19445_),
    .B(\count_cycle[32] ),
    .C(_19446_),
    .Y(_19447_));
 sky130_fd_sc_hd__nor2_4 _22476_ (.A(_19422_),
    .B(_19447_),
    .Y(_19448_));
 sky130_vsdinv _22477_ (.A(\count_cycle[34] ),
    .Y(_19449_));
 sky130_vsdinv _22478_ (.A(\count_cycle[35] ),
    .Y(_19450_));
 sky130_fd_sc_hd__nor2_2 _22479_ (.A(_19449_),
    .B(_19450_),
    .Y(_19451_));
 sky130_vsdinv _22480_ (.A(\count_cycle[36] ),
    .Y(_19452_));
 sky130_vsdinv _22481_ (.A(\count_cycle[37] ),
    .Y(_19453_));
 sky130_fd_sc_hd__nor2_2 _22482_ (.A(_19452_),
    .B(_19453_),
    .Y(_19454_));
 sky130_fd_sc_hd__nand3_4 _22483_ (.A(_19448_),
    .B(_19451_),
    .C(_19454_),
    .Y(_19455_));
 sky130_fd_sc_hd__nor3_4 _22484_ (.A(_19413_),
    .B(_19418_),
    .C(_19455_),
    .Y(_19456_));
 sky130_vsdinv _22485_ (.A(\count_cycle[47] ),
    .Y(_19457_));
 sky130_vsdinv _22486_ (.A(\count_cycle[45] ),
    .Y(_19458_));
 sky130_vsdinv _22487_ (.A(\count_cycle[46] ),
    .Y(_19459_));
 sky130_fd_sc_hd__or3b_4 _22488_ (.A(_19458_),
    .B(_19459_),
    .C_N(\count_cycle[44] ),
    .X(_19460_));
 sky130_fd_sc_hd__nor2_4 _22489_ (.A(_19457_),
    .B(_19460_),
    .Y(_19461_));
 sky130_fd_sc_hd__and3_1 _22490_ (.A(\count_cycle[48] ),
    .B(\count_cycle[49] ),
    .C(\count_cycle[50] ),
    .X(_19462_));
 sky130_fd_sc_hd__nand3_4 _22491_ (.A(_19456_),
    .B(_19461_),
    .C(_19462_),
    .Y(_19463_));
 sky130_fd_sc_hd__nor3_4 _22492_ (.A(_19404_),
    .B(_19409_),
    .C(_19463_),
    .Y(_19464_));
 sky130_fd_sc_hd__clkbuf_2 _22493_ (.A(_19464_),
    .X(_19465_));
 sky130_fd_sc_hd__and3_1 _22494_ (.A(\count_cycle[57] ),
    .B(\count_cycle[58] ),
    .C(\count_cycle[59] ),
    .X(_19466_));
 sky130_fd_sc_hd__clkbuf_2 _22495_ (.A(_19466_),
    .X(_19467_));
 sky130_fd_sc_hd__and3_1 _22496_ (.A(\count_cycle[60] ),
    .B(\count_cycle[61] ),
    .C(\count_cycle[62] ),
    .X(_19468_));
 sky130_fd_sc_hd__a41o_1 _22497_ (.A1(_19465_),
    .A2(\count_cycle[63] ),
    .A3(_19467_),
    .A4(_19468_),
    .B1(_19158_),
    .X(_19469_));
 sky130_fd_sc_hd__a31o_1 _22498_ (.A1(_19464_),
    .A2(_19466_),
    .A3(_19468_),
    .B1(\count_cycle[63] ),
    .X(_19470_));
 sky130_fd_sc_hd__nor2b_1 _22499_ (.A(_19469_),
    .B_N(_19470_),
    .Y(_03794_));
 sky130_fd_sc_hd__a31o_1 _22500_ (.A1(_19465_),
    .A2(_19467_),
    .A3(_19468_),
    .B1(_19158_),
    .X(_19471_));
 sky130_fd_sc_hd__clkbuf_2 _22501_ (.A(\count_cycle[60] ),
    .X(_19472_));
 sky130_fd_sc_hd__a41o_1 _22502_ (.A1(_19464_),
    .A2(_19472_),
    .A3(\count_cycle[61] ),
    .A4(_19466_),
    .B1(\count_cycle[62] ),
    .X(_19473_));
 sky130_fd_sc_hd__nor2b_1 _22503_ (.A(_19471_),
    .B_N(_19473_),
    .Y(_03793_));
 sky130_fd_sc_hd__a41o_1 _22504_ (.A1(_19465_),
    .A2(_19472_),
    .A3(\count_cycle[61] ),
    .A4(_19467_),
    .B1(_19158_),
    .X(_19474_));
 sky130_fd_sc_hd__a31o_1 _22505_ (.A1(_19464_),
    .A2(_19472_),
    .A3(_19466_),
    .B1(\count_cycle[61] ),
    .X(_19475_));
 sky130_fd_sc_hd__nor2b_1 _22506_ (.A(_19474_),
    .B_N(_19475_),
    .Y(_03792_));
 sky130_fd_sc_hd__buf_2 _22507_ (.A(_19464_),
    .X(_19476_));
 sky130_fd_sc_hd__a21oi_1 _22508_ (.A1(_19476_),
    .A2(_19467_),
    .B1(_19472_),
    .Y(_19477_));
 sky130_fd_sc_hd__a31o_1 _22509_ (.A1(_19465_),
    .A2(_19472_),
    .A3(_19467_),
    .B1(_19158_),
    .X(_19478_));
 sky130_fd_sc_hd__nor2_1 _22510_ (.A(_19477_),
    .B(_19478_),
    .Y(_03791_));
 sky130_fd_sc_hd__nand2_1 _22511_ (.A(\count_cycle[57] ),
    .B(\count_cycle[58] ),
    .Y(_19479_));
 sky130_vsdinv _22512_ (.A(_19479_),
    .Y(_19480_));
 sky130_fd_sc_hd__a21oi_1 _22513_ (.A1(_19465_),
    .A2(_19480_),
    .B1(\count_cycle[59] ),
    .Y(_19481_));
 sky130_fd_sc_hd__a211oi_2 _22514_ (.A1(_19476_),
    .A2(_19467_),
    .B1(_18794_),
    .C1(_19481_),
    .Y(_03790_));
 sky130_fd_sc_hd__a21oi_1 _22515_ (.A1(_19465_),
    .A2(\count_cycle[57] ),
    .B1(\count_cycle[58] ),
    .Y(_19482_));
 sky130_fd_sc_hd__a211oi_2 _22516_ (.A1(_19476_),
    .A2(_19480_),
    .B1(_18794_),
    .C1(_19482_),
    .Y(_03789_));
 sky130_fd_sc_hd__a21oi_1 _22517_ (.A1(_19476_),
    .A2(\count_cycle[57] ),
    .B1(_18757_),
    .Y(_19483_));
 sky130_fd_sc_hd__o21a_1 _22518_ (.A1(\count_cycle[57] ),
    .A2(_19476_),
    .B1(_19483_),
    .X(_03788_));
 sky130_fd_sc_hd__buf_2 _22519_ (.A(_19463_),
    .X(_19484_));
 sky130_fd_sc_hd__nor2_1 _22520_ (.A(_19409_),
    .B(_19484_),
    .Y(_19485_));
 sky130_fd_sc_hd__o21ai_1 _22521_ (.A1(\count_cycle[56] ),
    .A2(_19485_),
    .B1(_19175_),
    .Y(_19486_));
 sky130_fd_sc_hd__nor2_1 _22522_ (.A(_19476_),
    .B(_19486_),
    .Y(_03787_));
 sky130_fd_sc_hd__nor3_4 _22523_ (.A(_19406_),
    .B(_19407_),
    .C(_19484_),
    .Y(_19487_));
 sky130_fd_sc_hd__a31o_1 _22524_ (.A1(_19487_),
    .A2(\count_cycle[53] ),
    .A3(\count_cycle[54] ),
    .B1(\count_cycle[55] ),
    .X(_19488_));
 sky130_fd_sc_hd__o211a_1 _22525_ (.A1(_19484_),
    .A2(_19409_),
    .B1(_19195_),
    .C1(_19488_),
    .X(_03786_));
 sky130_vsdinv _22526_ (.A(_19487_),
    .Y(_19489_));
 sky130_fd_sc_hd__nor2_1 _22527_ (.A(_19408_),
    .B(_19489_),
    .Y(_19490_));
 sky130_fd_sc_hd__a31o_1 _22528_ (.A1(_19487_),
    .A2(\count_cycle[53] ),
    .A3(\count_cycle[54] ),
    .B1(_18793_),
    .X(_19491_));
 sky130_fd_sc_hd__o21ba_1 _22529_ (.A1(\count_cycle[54] ),
    .A2(_19490_),
    .B1_N(_19491_),
    .X(_03785_));
 sky130_fd_sc_hd__nor2_1 _22530_ (.A(\count_cycle[53] ),
    .B(_19487_),
    .Y(_19492_));
 sky130_fd_sc_hd__nor3_1 _22531_ (.A(_19179_),
    .B(_19492_),
    .C(_19490_),
    .Y(_03784_));
 sky130_fd_sc_hd__or2_1 _22532_ (.A(_19406_),
    .B(_19484_),
    .X(_19493_));
 sky130_fd_sc_hd__nand2_1 _22533_ (.A(_19493_),
    .B(_19407_),
    .Y(_19494_));
 sky130_fd_sc_hd__and3_1 _22534_ (.A(_19494_),
    .B(_19489_),
    .C(_19195_),
    .X(_03783_));
 sky130_fd_sc_hd__nand2_1 _22535_ (.A(_19484_),
    .B(_19406_),
    .Y(_19495_));
 sky130_fd_sc_hd__and3_1 _22536_ (.A(_19493_),
    .B(_19308_),
    .C(_19495_),
    .X(_03782_));
 sky130_vsdinv _22537_ (.A(\count_cycle[49] ),
    .Y(_19496_));
 sky130_fd_sc_hd__nand3_2 _22538_ (.A(_19456_),
    .B(\count_cycle[48] ),
    .C(_19461_),
    .Y(_19497_));
 sky130_fd_sc_hd__nor2_1 _22539_ (.A(_19496_),
    .B(_19497_),
    .Y(_19498_));
 sky130_fd_sc_hd__or2_1 _22540_ (.A(\count_cycle[50] ),
    .B(_19498_),
    .X(_19499_));
 sky130_fd_sc_hd__clkbuf_2 _22541_ (.A(_19244_),
    .X(_19500_));
 sky130_fd_sc_hd__and3_1 _22542_ (.A(_19499_),
    .B(_19500_),
    .C(_19484_),
    .X(_03781_));
 sky130_fd_sc_hd__or2_1 _22543_ (.A(_19252_),
    .B(_19498_),
    .X(_19501_));
 sky130_fd_sc_hd__a21oi_1 _22544_ (.A1(_19496_),
    .A2(_19497_),
    .B1(_19501_),
    .Y(_03780_));
 sky130_fd_sc_hd__and2_1 _22545_ (.A(_19456_),
    .B(_19461_),
    .X(_19502_));
 sky130_fd_sc_hd__or2_1 _22546_ (.A(\count_cycle[48] ),
    .B(_19502_),
    .X(_19503_));
 sky130_fd_sc_hd__and3_1 _22547_ (.A(_19503_),
    .B(_19500_),
    .C(_19497_),
    .X(_03779_));
 sky130_vsdinv _22548_ (.A(_19456_),
    .Y(_19504_));
 sky130_fd_sc_hd__or2_1 _22549_ (.A(_19460_),
    .B(_19504_),
    .X(_19505_));
 sky130_fd_sc_hd__clkbuf_4 _22550_ (.A(_18557_),
    .X(_19506_));
 sky130_fd_sc_hd__or2_1 _22551_ (.A(_19506_),
    .B(_19502_),
    .X(_19507_));
 sky130_fd_sc_hd__a21oi_1 _22552_ (.A1(_19505_),
    .A2(_19457_),
    .B1(_19507_),
    .Y(_03778_));
 sky130_fd_sc_hd__nand2_1 _22553_ (.A(_19456_),
    .B(\count_cycle[44] ),
    .Y(_19508_));
 sky130_fd_sc_hd__or2_1 _22554_ (.A(_19458_),
    .B(_19508_),
    .X(_19509_));
 sky130_fd_sc_hd__nand2_1 _22555_ (.A(_19509_),
    .B(_19459_),
    .Y(_19510_));
 sky130_fd_sc_hd__and3_1 _22556_ (.A(_19510_),
    .B(_19500_),
    .C(_19505_),
    .X(_03777_));
 sky130_fd_sc_hd__nand2_1 _22557_ (.A(_19508_),
    .B(_19458_),
    .Y(_19511_));
 sky130_fd_sc_hd__and3_1 _22558_ (.A(_19509_),
    .B(_19500_),
    .C(_19511_),
    .X(_03776_));
 sky130_fd_sc_hd__or2_1 _22559_ (.A(\count_cycle[44] ),
    .B(_19456_),
    .X(_19512_));
 sky130_fd_sc_hd__and3_1 _22560_ (.A(_19512_),
    .B(_19500_),
    .C(_19508_),
    .X(_03775_));
 sky130_fd_sc_hd__nor3_4 _22561_ (.A(_19414_),
    .B(_19413_),
    .C(_19455_),
    .Y(_19513_));
 sky130_fd_sc_hd__nand2_1 _22562_ (.A(_19513_),
    .B(\count_cycle[41] ),
    .Y(_19514_));
 sky130_fd_sc_hd__or2_1 _22563_ (.A(_19416_),
    .B(_19514_),
    .X(_19515_));
 sky130_fd_sc_hd__nand2_1 _22564_ (.A(_19515_),
    .B(_19417_),
    .Y(_19516_));
 sky130_fd_sc_hd__and3_1 _22565_ (.A(_19516_),
    .B(_19500_),
    .C(_19504_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_2 _22566_ (.A(_19244_),
    .X(_19517_));
 sky130_fd_sc_hd__nand2_1 _22567_ (.A(_19514_),
    .B(_19416_),
    .Y(_19518_));
 sky130_fd_sc_hd__and3_1 _22568_ (.A(_19515_),
    .B(_19517_),
    .C(_19518_),
    .X(_03773_));
 sky130_fd_sc_hd__or2_1 _22569_ (.A(\count_cycle[41] ),
    .B(_19513_),
    .X(_19519_));
 sky130_fd_sc_hd__and3_1 _22570_ (.A(_19519_),
    .B(_19517_),
    .C(_19514_),
    .X(_03772_));
 sky130_fd_sc_hd__or2_1 _22571_ (.A(_19413_),
    .B(_19455_),
    .X(_19520_));
 sky130_fd_sc_hd__or2_1 _22572_ (.A(_19506_),
    .B(_19513_),
    .X(_19521_));
 sky130_fd_sc_hd__a21oi_1 _22573_ (.A1(_19414_),
    .A2(_19520_),
    .B1(_19521_),
    .Y(_03771_));
 sky130_fd_sc_hd__or2_1 _22574_ (.A(_19410_),
    .B(_19455_),
    .X(_19522_));
 sky130_fd_sc_hd__nand2_1 _22575_ (.A(_19522_),
    .B(_19411_),
    .Y(_19523_));
 sky130_fd_sc_hd__and3_1 _22576_ (.A(_19523_),
    .B(_19517_),
    .C(_19520_),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_1 _22577_ (.A(_19455_),
    .B(_19410_),
    .Y(_19524_));
 sky130_fd_sc_hd__and3_1 _22578_ (.A(_19522_),
    .B(_19517_),
    .C(_19524_),
    .X(_03769_));
 sky130_fd_sc_hd__nand2_1 _22579_ (.A(_19448_),
    .B(_19451_),
    .Y(_19525_));
 sky130_fd_sc_hd__or2_1 _22580_ (.A(_19452_),
    .B(_19525_),
    .X(_19526_));
 sky130_fd_sc_hd__nand2_1 _22581_ (.A(_19526_),
    .B(_19453_),
    .Y(_19527_));
 sky130_fd_sc_hd__and3_1 _22582_ (.A(_19527_),
    .B(_19517_),
    .C(_19455_),
    .X(_03768_));
 sky130_fd_sc_hd__nand2_1 _22583_ (.A(_19525_),
    .B(_19452_),
    .Y(_19528_));
 sky130_fd_sc_hd__and3_1 _22584_ (.A(_19526_),
    .B(_19517_),
    .C(_19528_),
    .X(_03767_));
 sky130_fd_sc_hd__nand2_1 _22585_ (.A(_19448_),
    .B(\count_cycle[34] ),
    .Y(_19529_));
 sky130_fd_sc_hd__nand2_1 _22586_ (.A(_19529_),
    .B(_19450_),
    .Y(_19530_));
 sky130_fd_sc_hd__buf_1 _22587_ (.A(_19188_),
    .X(_19531_));
 sky130_fd_sc_hd__and3_1 _22588_ (.A(_19530_),
    .B(_19531_),
    .C(_19525_),
    .X(_03766_));
 sky130_vsdinv _22589_ (.A(_19448_),
    .Y(_19532_));
 sky130_fd_sc_hd__nand2_1 _22590_ (.A(_19532_),
    .B(_19449_),
    .Y(_19533_));
 sky130_fd_sc_hd__and3_1 _22591_ (.A(_19533_),
    .B(_19531_),
    .C(_19529_),
    .X(_03765_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(_19420_),
    .B(_19447_),
    .Y(_19534_));
 sky130_vsdinv _22593_ (.A(_19534_),
    .Y(_19535_));
 sky130_fd_sc_hd__nand2_1 _22594_ (.A(_19535_),
    .B(_19419_),
    .Y(_19536_));
 sky130_fd_sc_hd__and3_1 _22595_ (.A(_19536_),
    .B(_19531_),
    .C(_19532_),
    .X(_03764_));
 sky130_fd_sc_hd__nand2_1 _22596_ (.A(_19445_),
    .B(_19446_),
    .Y(_19537_));
 sky130_fd_sc_hd__or2_1 _22597_ (.A(_19420_),
    .B(_19537_),
    .X(_19538_));
 sky130_vsdinv _22598_ (.A(\count_cycle[32] ),
    .Y(_19539_));
 sky130_fd_sc_hd__nand2_1 _22599_ (.A(_19538_),
    .B(_19539_),
    .Y(_19540_));
 sky130_fd_sc_hd__and3_1 _22600_ (.A(_19540_),
    .B(_19531_),
    .C(_19535_),
    .X(_03763_));
 sky130_fd_sc_hd__or2_1 _22601_ (.A(_02028_),
    .B(_19537_),
    .X(_19541_));
 sky130_fd_sc_hd__or2_1 _22602_ (.A(_02037_),
    .B(_19541_),
    .X(_19542_));
 sky130_fd_sc_hd__or2_1 _22603_ (.A(_02046_),
    .B(_19542_),
    .X(_19543_));
 sky130_fd_sc_hd__nand2_1 _22604_ (.A(_19543_),
    .B(_02055_),
    .Y(_19544_));
 sky130_fd_sc_hd__and3_1 _22605_ (.A(_19544_),
    .B(_19531_),
    .C(_19538_),
    .X(_03762_));
 sky130_fd_sc_hd__nand2_1 _22606_ (.A(_19542_),
    .B(_02046_),
    .Y(_19545_));
 sky130_fd_sc_hd__and3_1 _22607_ (.A(_19543_),
    .B(_19531_),
    .C(_19545_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_2 _22608_ (.A(_19188_),
    .X(_19546_));
 sky130_fd_sc_hd__nand2_1 _22609_ (.A(_19541_),
    .B(_02037_),
    .Y(_19547_));
 sky130_fd_sc_hd__and3_1 _22610_ (.A(_19542_),
    .B(_19546_),
    .C(_19547_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_1 _22611_ (.A(_19537_),
    .B(_02028_),
    .Y(_19548_));
 sky130_fd_sc_hd__and3_1 _22612_ (.A(_19541_),
    .B(_19546_),
    .C(_19548_),
    .X(_03759_));
 sky130_fd_sc_hd__nand2_1 _22613_ (.A(_19445_),
    .B(\count_cycle[26] ),
    .Y(_19549_));
 sky130_fd_sc_hd__nand2_1 _22614_ (.A(_19549_),
    .B(_02019_),
    .Y(_19550_));
 sky130_fd_sc_hd__and3_1 _22615_ (.A(_19550_),
    .B(_19546_),
    .C(_19537_),
    .X(_03758_));
 sky130_fd_sc_hd__or2_1 _22616_ (.A(\count_cycle[26] ),
    .B(_19445_),
    .X(_19551_));
 sky130_fd_sc_hd__and3_1 _22617_ (.A(_19551_),
    .B(_19546_),
    .C(_19549_),
    .X(_03757_));
 sky130_fd_sc_hd__nand2_1 _22618_ (.A(_19443_),
    .B(\count_cycle[23] ),
    .Y(_19552_));
 sky130_fd_sc_hd__nor2_1 _22619_ (.A(_01992_),
    .B(_19552_),
    .Y(_19553_));
 sky130_fd_sc_hd__nor2_1 _22620_ (.A(_18843_),
    .B(_19445_),
    .Y(_19554_));
 sky130_fd_sc_hd__o21a_1 _22621_ (.A1(\count_cycle[25] ),
    .A2(_19553_),
    .B1(_19554_),
    .X(_03756_));
 sky130_fd_sc_hd__or2_1 _22622_ (.A(_19506_),
    .B(_19553_),
    .X(_19555_));
 sky130_fd_sc_hd__a21oi_1 _22623_ (.A1(_01992_),
    .A2(_19552_),
    .B1(_19555_),
    .Y(_03755_));
 sky130_vsdinv _22624_ (.A(_19443_),
    .Y(_19556_));
 sky130_fd_sc_hd__nand2_1 _22625_ (.A(_19556_),
    .B(_01983_),
    .Y(_19557_));
 sky130_fd_sc_hd__and3_1 _22626_ (.A(_19557_),
    .B(_19546_),
    .C(_19552_),
    .X(_03754_));
 sky130_fd_sc_hd__nand2_1 _22627_ (.A(_19442_),
    .B(_01974_),
    .Y(_19558_));
 sky130_fd_sc_hd__and3_1 _22628_ (.A(_19556_),
    .B(_19546_),
    .C(_19558_),
    .X(_03753_));
 sky130_vsdinv _22629_ (.A(_19441_),
    .Y(_19559_));
 sky130_fd_sc_hd__inv_2 _22630_ (.A(\count_cycle[21] ),
    .Y(_01965_));
 sky130_fd_sc_hd__nand2_1 _22631_ (.A(_19559_),
    .B(_01965_),
    .Y(_19560_));
 sky130_fd_sc_hd__clkbuf_2 _22632_ (.A(_19188_),
    .X(_19561_));
 sky130_fd_sc_hd__and3_1 _22633_ (.A(_19560_),
    .B(_19561_),
    .C(_19442_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _22634_ (.A(_19440_),
    .B(_01956_),
    .Y(_19562_));
 sky130_fd_sc_hd__and3_1 _22635_ (.A(_19559_),
    .B(_19561_),
    .C(_19562_),
    .X(_03751_));
 sky130_fd_sc_hd__or2_1 _22636_ (.A(\count_cycle[19] ),
    .B(_19439_),
    .X(_19563_));
 sky130_fd_sc_hd__and3_1 _22637_ (.A(_19563_),
    .B(_19561_),
    .C(_19440_),
    .X(_03750_));
 sky130_fd_sc_hd__or2_1 _22638_ (.A(_19506_),
    .B(_19439_),
    .X(_19564_));
 sky130_fd_sc_hd__a21oi_1 _22639_ (.A1(_01938_),
    .A2(_19438_),
    .B1(_19564_),
    .Y(_03749_));
 sky130_vsdinv _22640_ (.A(_19437_),
    .Y(_19565_));
 sky130_fd_sc_hd__inv_2 _22641_ (.A(\count_cycle[17] ),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_1 _22642_ (.A(_19565_),
    .B(_01929_),
    .Y(_19566_));
 sky130_fd_sc_hd__and3_1 _22643_ (.A(_19566_),
    .B(_19561_),
    .C(_19438_),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_1 _22644_ (.A(_19436_),
    .B(_01920_),
    .Y(_19567_));
 sky130_fd_sc_hd__and3_1 _22645_ (.A(_19565_),
    .B(_19561_),
    .C(_19567_),
    .X(_03747_));
 sky130_fd_sc_hd__nand2_1 _22646_ (.A(_19435_),
    .B(_01911_),
    .Y(_19568_));
 sky130_fd_sc_hd__and3_1 _22647_ (.A(_19436_),
    .B(_19561_),
    .C(_19568_),
    .X(_03746_));
 sky130_fd_sc_hd__or2_1 _22648_ (.A(\count_cycle[14] ),
    .B(_19434_),
    .X(_19569_));
 sky130_fd_sc_hd__clkbuf_2 _22649_ (.A(_19188_),
    .X(_19570_));
 sky130_fd_sc_hd__and3_1 _22650_ (.A(_19569_),
    .B(_19570_),
    .C(_19435_),
    .X(_03745_));
 sky130_fd_sc_hd__or2_1 _22651_ (.A(_19506_),
    .B(_19434_),
    .X(_19571_));
 sky130_fd_sc_hd__a21oi_1 _22652_ (.A1(_01885_),
    .A2(_19433_),
    .B1(_19571_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _22653_ (.A(_19432_),
    .B(_01872_),
    .Y(_19572_));
 sky130_fd_sc_hd__and3_1 _22654_ (.A(_19433_),
    .B(_19570_),
    .C(_19572_),
    .X(_03743_));
 sky130_vsdinv _22655_ (.A(_19431_),
    .Y(_19573_));
 sky130_fd_sc_hd__inv_2 _22656_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _22657_ (.A(_19573_),
    .B(_01859_),
    .Y(_19574_));
 sky130_fd_sc_hd__and3_1 _22658_ (.A(_19574_),
    .B(_19570_),
    .C(_19432_),
    .X(_03742_));
 sky130_fd_sc_hd__nand2_1 _22659_ (.A(_19430_),
    .B(_01846_),
    .Y(_19575_));
 sky130_fd_sc_hd__and3_1 _22660_ (.A(_19573_),
    .B(_19570_),
    .C(_19575_),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_1 _22661_ (.A(_19429_),
    .B(_01833_),
    .Y(_19576_));
 sky130_fd_sc_hd__and3_1 _22662_ (.A(_19430_),
    .B(_19570_),
    .C(_19576_),
    .X(_03740_));
 sky130_fd_sc_hd__or2_1 _22663_ (.A(_01806_),
    .B(_19428_),
    .X(_19577_));
 sky130_fd_sc_hd__nand2_1 _22664_ (.A(_19577_),
    .B(_01820_),
    .Y(_19578_));
 sky130_fd_sc_hd__and3_1 _22665_ (.A(_19578_),
    .B(_19429_),
    .C(_19189_),
    .X(_03739_));
 sky130_fd_sc_hd__nand2_1 _22666_ (.A(_19428_),
    .B(_01806_),
    .Y(_19579_));
 sky130_fd_sc_hd__and3_1 _22667_ (.A(_19577_),
    .B(_19570_),
    .C(_19579_),
    .X(_03738_));
 sky130_vsdinv _22668_ (.A(_19427_),
    .Y(_19580_));
 sky130_fd_sc_hd__inv_2 _22669_ (.A(\count_cycle[6] ),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _22670_ (.A(_19580_),
    .B(_01793_),
    .Y(_19581_));
 sky130_fd_sc_hd__buf_1 _22671_ (.A(_19188_),
    .X(_19582_));
 sky130_fd_sc_hd__and3_1 _22672_ (.A(_19581_),
    .B(_19582_),
    .C(_19428_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_1 _22673_ (.A(_19426_),
    .B(_01780_),
    .Y(_19583_));
 sky130_fd_sc_hd__and3_1 _22674_ (.A(_19580_),
    .B(_19582_),
    .C(_19583_),
    .X(_03736_));
 sky130_vsdinv _22675_ (.A(_19425_),
    .Y(_19584_));
 sky130_fd_sc_hd__inv_2 _22676_ (.A(\count_cycle[4] ),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _22677_ (.A(_19584_),
    .B(_01767_),
    .Y(_19585_));
 sky130_fd_sc_hd__and3_1 _22678_ (.A(_19585_),
    .B(_19582_),
    .C(_19426_),
    .X(_03735_));
 sky130_fd_sc_hd__nand2_1 _22679_ (.A(_19424_),
    .B(_01754_),
    .Y(_19586_));
 sky130_fd_sc_hd__and3_1 _22680_ (.A(_19584_),
    .B(_19582_),
    .C(_19586_),
    .X(_03734_));
 sky130_fd_sc_hd__nand2_1 _22681_ (.A(_01741_),
    .B(_19423_),
    .Y(_19587_));
 sky130_fd_sc_hd__and3_1 _22682_ (.A(_19424_),
    .B(_19582_),
    .C(_19587_),
    .X(_03733_));
 sky130_fd_sc_hd__inv_2 _22683_ (.A(\count_cycle[0] ),
    .Y(_02559_));
 sky130_fd_sc_hd__inv_2 _22684_ (.A(\count_cycle[1] ),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_1 _22685_ (.A(_02559_),
    .B(_01728_),
    .Y(_19588_));
 sky130_fd_sc_hd__and3_1 _22686_ (.A(_19588_),
    .B(_19582_),
    .C(_19423_),
    .X(_03732_));
 sky130_fd_sc_hd__nor2_1 _22687_ (.A(\count_cycle[0] ),
    .B(_18867_),
    .Y(_03731_));
 sky130_fd_sc_hd__nor2_1 _22688_ (.A(_18758_),
    .B(_18962_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _22689_ (.A(_18758_),
    .B(_18676_),
    .Y(_03729_));
 sky130_vsdinv _22690_ (.A(_18689_),
    .Y(_03728_));
 sky130_fd_sc_hd__clkbuf_2 _22691_ (.A(\cpuregs_wrdata[31] ),
    .X(_19589_));
 sky130_vsdinv _22692_ (.A(\latched_rd[1] ),
    .Y(_19590_));
 sky130_vsdinv _22693_ (.A(\latched_rd[0] ),
    .Y(_19591_));
 sky130_fd_sc_hd__nand2_2 _22694_ (.A(_19591_),
    .B(_19590_),
    .Y(_19592_));
 sky130_fd_sc_hd__nor2_1 _22695_ (.A(\latched_rd[4] ),
    .B(\latched_rd[2] ),
    .Y(_19593_));
 sky130_vsdinv _22696_ (.A(\latched_rd[3] ),
    .Y(_19594_));
 sky130_fd_sc_hd__nand2_2 _22697_ (.A(_19593_),
    .B(_19594_),
    .Y(_19595_));
 sky130_vsdinv _22698_ (.A(_18656_),
    .Y(_19596_));
 sky130_fd_sc_hd__nor2_4 _22699_ (.A(_18531_),
    .B(_18720_),
    .Y(_19597_));
 sky130_fd_sc_hd__o31a_4 _22700_ (.A1(latched_branch),
    .A2(net511),
    .A3(_19596_),
    .B1(_19597_),
    .X(_19598_));
 sky130_fd_sc_hd__o21ai_4 _22701_ (.A1(_19592_),
    .A2(_19595_),
    .B1(_19598_),
    .Y(_19599_));
 sky130_fd_sc_hd__or2_2 _22702_ (.A(_19590_),
    .B(_19599_),
    .X(_19600_));
 sky130_fd_sc_hd__nor2_4 _22703_ (.A(\latched_rd[0] ),
    .B(_19600_),
    .Y(_19601_));
 sky130_vsdinv _22704_ (.A(\latched_rd[4] ),
    .Y(_19602_));
 sky130_fd_sc_hd__and3_1 _22705_ (.A(_19602_),
    .B(_19594_),
    .C(\latched_rd[2] ),
    .X(_19603_));
 sky130_fd_sc_hd__nand2_1 _22706_ (.A(_19601_),
    .B(_19603_),
    .Y(_19604_));
 sky130_fd_sc_hd__buf_6 _22707_ (.A(_19604_),
    .X(_19605_));
 sky130_fd_sc_hd__clkbuf_4 _22708_ (.A(_19605_),
    .X(_19606_));
 sky130_fd_sc_hd__mux2_1 _22709_ (.A0(_19589_),
    .A1(\cpuregs[6][31] ),
    .S(_19606_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_2 _22710_ (.A(\cpuregs_wrdata[30] ),
    .X(_19607_));
 sky130_fd_sc_hd__mux2_1 _22711_ (.A0(_19607_),
    .A1(\cpuregs[6][30] ),
    .S(_19606_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_2 _22712_ (.A(\cpuregs_wrdata[29] ),
    .X(_19608_));
 sky130_fd_sc_hd__mux2_1 _22713_ (.A0(_19608_),
    .A1(\cpuregs[6][29] ),
    .S(_19606_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_2 _22714_ (.A(\cpuregs_wrdata[28] ),
    .X(_19609_));
 sky130_fd_sc_hd__mux2_1 _22715_ (.A0(_19609_),
    .A1(\cpuregs[6][28] ),
    .S(_19606_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_2 _22716_ (.A(\cpuregs_wrdata[27] ),
    .X(_19610_));
 sky130_fd_sc_hd__mux2_1 _22717_ (.A0(_19610_),
    .A1(\cpuregs[6][27] ),
    .S(_19606_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_2 _22718_ (.A(\cpuregs_wrdata[26] ),
    .X(_19611_));
 sky130_fd_sc_hd__mux2_1 _22719_ (.A0(_19611_),
    .A1(\cpuregs[6][26] ),
    .S(_19606_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_2 _22720_ (.A(\cpuregs_wrdata[25] ),
    .X(_19612_));
 sky130_fd_sc_hd__clkbuf_4 _22721_ (.A(_19605_),
    .X(_19613_));
 sky130_fd_sc_hd__mux2_1 _22722_ (.A0(_19612_),
    .A1(\cpuregs[6][25] ),
    .S(_19613_),
    .X(_03721_));
 sky130_fd_sc_hd__buf_1 _22723_ (.A(\cpuregs_wrdata[24] ),
    .X(_19614_));
 sky130_fd_sc_hd__mux2_1 _22724_ (.A0(_19614_),
    .A1(\cpuregs[6][24] ),
    .S(_19613_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_2 _22725_ (.A(\cpuregs_wrdata[23] ),
    .X(_19615_));
 sky130_fd_sc_hd__mux2_1 _22726_ (.A0(_19615_),
    .A1(\cpuregs[6][23] ),
    .S(_19613_),
    .X(_03719_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22727_ (.A(\cpuregs_wrdata[22] ),
    .X(_19616_));
 sky130_fd_sc_hd__mux2_1 _22728_ (.A0(_19616_),
    .A1(\cpuregs[6][22] ),
    .S(_19613_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_2 _22729_ (.A(\cpuregs_wrdata[21] ),
    .X(_19617_));
 sky130_fd_sc_hd__mux2_1 _22730_ (.A0(_19617_),
    .A1(\cpuregs[6][21] ),
    .S(_19613_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_2 _22731_ (.A(\cpuregs_wrdata[20] ),
    .X(_19618_));
 sky130_fd_sc_hd__mux2_1 _22732_ (.A0(_19618_),
    .A1(\cpuregs[6][20] ),
    .S(_19613_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_2 _22733_ (.A(\cpuregs_wrdata[19] ),
    .X(_19619_));
 sky130_fd_sc_hd__buf_2 _22734_ (.A(_19605_),
    .X(_19620_));
 sky130_fd_sc_hd__mux2_1 _22735_ (.A0(_19619_),
    .A1(\cpuregs[6][19] ),
    .S(_19620_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_2 _22736_ (.A(\cpuregs_wrdata[18] ),
    .X(_19621_));
 sky130_fd_sc_hd__mux2_1 _22737_ (.A0(_19621_),
    .A1(\cpuregs[6][18] ),
    .S(_19620_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_2 _22738_ (.A(\cpuregs_wrdata[17] ),
    .X(_19622_));
 sky130_fd_sc_hd__mux2_1 _22739_ (.A0(_19622_),
    .A1(\cpuregs[6][17] ),
    .S(_19620_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_2 _22740_ (.A(\cpuregs_wrdata[16] ),
    .X(_19623_));
 sky130_fd_sc_hd__mux2_1 _22741_ (.A0(_19623_),
    .A1(\cpuregs[6][16] ),
    .S(_19620_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_2 _22742_ (.A(\cpuregs_wrdata[15] ),
    .X(_19624_));
 sky130_fd_sc_hd__mux2_1 _22743_ (.A0(_19624_),
    .A1(\cpuregs[6][15] ),
    .S(_19620_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_2 _22744_ (.A(\cpuregs_wrdata[14] ),
    .X(_19625_));
 sky130_fd_sc_hd__mux2_1 _22745_ (.A0(_19625_),
    .A1(\cpuregs[6][14] ),
    .S(_19620_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_2 _22746_ (.A(\cpuregs_wrdata[13] ),
    .X(_19626_));
 sky130_fd_sc_hd__clkbuf_4 _22747_ (.A(_19605_),
    .X(_19627_));
 sky130_fd_sc_hd__mux2_1 _22748_ (.A0(_19626_),
    .A1(\cpuregs[6][13] ),
    .S(_19627_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_2 _22749_ (.A(\cpuregs_wrdata[12] ),
    .X(_19628_));
 sky130_fd_sc_hd__mux2_1 _22750_ (.A0(_19628_),
    .A1(\cpuregs[6][12] ),
    .S(_19627_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_2 _22751_ (.A(\cpuregs_wrdata[11] ),
    .X(_19629_));
 sky130_fd_sc_hd__mux2_1 _22752_ (.A0(_19629_),
    .A1(\cpuregs[6][11] ),
    .S(_19627_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_2 _22753_ (.A(\cpuregs_wrdata[10] ),
    .X(_19630_));
 sky130_fd_sc_hd__mux2_1 _22754_ (.A0(_19630_),
    .A1(\cpuregs[6][10] ),
    .S(_19627_),
    .X(_03706_));
 sky130_fd_sc_hd__buf_1 _22755_ (.A(\cpuregs_wrdata[9] ),
    .X(_19631_));
 sky130_fd_sc_hd__mux2_1 _22756_ (.A0(_19631_),
    .A1(\cpuregs[6][9] ),
    .S(_19627_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_2 _22757_ (.A(\cpuregs_wrdata[8] ),
    .X(_19632_));
 sky130_fd_sc_hd__mux2_1 _22758_ (.A0(_19632_),
    .A1(\cpuregs[6][8] ),
    .S(_19627_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_2 _22759_ (.A(\cpuregs_wrdata[7] ),
    .X(_19633_));
 sky130_fd_sc_hd__clkbuf_4 _22760_ (.A(_19604_),
    .X(_19634_));
 sky130_fd_sc_hd__mux2_1 _22761_ (.A0(_19633_),
    .A1(\cpuregs[6][7] ),
    .S(_19634_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_2 _22762_ (.A(\cpuregs_wrdata[6] ),
    .X(_19635_));
 sky130_fd_sc_hd__mux2_1 _22763_ (.A0(_19635_),
    .A1(\cpuregs[6][6] ),
    .S(_19634_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_2 _22764_ (.A(\cpuregs_wrdata[5] ),
    .X(_19636_));
 sky130_fd_sc_hd__mux2_1 _22765_ (.A0(_19636_),
    .A1(\cpuregs[6][5] ),
    .S(_19634_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_2 _22766_ (.A(\cpuregs_wrdata[4] ),
    .X(_19637_));
 sky130_fd_sc_hd__mux2_1 _22767_ (.A0(_19637_),
    .A1(\cpuregs[6][4] ),
    .S(_19634_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_2 _22768_ (.A(\cpuregs_wrdata[3] ),
    .X(_19638_));
 sky130_fd_sc_hd__mux2_1 _22769_ (.A0(_19638_),
    .A1(\cpuregs[6][3] ),
    .S(_19634_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_2 _22770_ (.A(\cpuregs_wrdata[2] ),
    .X(_19639_));
 sky130_fd_sc_hd__mux2_1 _22771_ (.A0(_19639_),
    .A1(\cpuregs[6][2] ),
    .S(_19634_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_2 _22772_ (.A(\cpuregs_wrdata[1] ),
    .X(_19640_));
 sky130_fd_sc_hd__mux2_1 _22773_ (.A0(_19640_),
    .A1(\cpuregs[6][1] ),
    .S(_19605_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_2 _22774_ (.A(\cpuregs_wrdata[0] ),
    .X(_19641_));
 sky130_fd_sc_hd__mux2_1 _22775_ (.A0(_19641_),
    .A1(\cpuregs[6][0] ),
    .S(_19605_),
    .X(_03696_));
 sky130_fd_sc_hd__nor3_4 _22776_ (.A(_19591_),
    .B(\latched_rd[1] ),
    .C(_19599_),
    .Y(_19642_));
 sky130_fd_sc_hd__nand2_1 _22777_ (.A(_19593_),
    .B(\latched_rd[3] ),
    .Y(_19643_));
 sky130_vsdinv _22778_ (.A(_19643_),
    .Y(_19644_));
 sky130_fd_sc_hd__nand2_1 _22779_ (.A(_19642_),
    .B(_19644_),
    .Y(_19645_));
 sky130_fd_sc_hd__buf_6 _22780_ (.A(_19645_),
    .X(_19646_));
 sky130_fd_sc_hd__clkbuf_4 _22781_ (.A(_19646_),
    .X(_19647_));
 sky130_fd_sc_hd__mux2_1 _22782_ (.A0(_19589_),
    .A1(\cpuregs[9][31] ),
    .S(_19647_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _22783_ (.A0(_19607_),
    .A1(\cpuregs[9][30] ),
    .S(_19647_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _22784_ (.A0(_19608_),
    .A1(\cpuregs[9][29] ),
    .S(_19647_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _22785_ (.A0(_19609_),
    .A1(\cpuregs[9][28] ),
    .S(_19647_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _22786_ (.A0(_19610_),
    .A1(\cpuregs[9][27] ),
    .S(_19647_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _22787_ (.A0(_19611_),
    .A1(\cpuregs[9][26] ),
    .S(_19647_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_4 _22788_ (.A(_19646_),
    .X(_19648_));
 sky130_fd_sc_hd__mux2_1 _22789_ (.A0(_19612_),
    .A1(\cpuregs[9][25] ),
    .S(_19648_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _22790_ (.A0(_19614_),
    .A1(\cpuregs[9][24] ),
    .S(_19648_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _22791_ (.A0(_19615_),
    .A1(\cpuregs[9][23] ),
    .S(_19648_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _22792_ (.A0(_19616_),
    .A1(\cpuregs[9][22] ),
    .S(_19648_),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_1 _22793_ (.A0(_19617_),
    .A1(\cpuregs[9][21] ),
    .S(_19648_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _22794_ (.A0(_19618_),
    .A1(\cpuregs[9][20] ),
    .S(_19648_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_4 _22795_ (.A(_19646_),
    .X(_19649_));
 sky130_fd_sc_hd__mux2_1 _22796_ (.A0(_19619_),
    .A1(\cpuregs[9][19] ),
    .S(_19649_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _22797_ (.A0(_19621_),
    .A1(\cpuregs[9][18] ),
    .S(_19649_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _22798_ (.A0(_19622_),
    .A1(\cpuregs[9][17] ),
    .S(_19649_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _22799_ (.A0(_19623_),
    .A1(\cpuregs[9][16] ),
    .S(_19649_),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _22800_ (.A0(_19624_),
    .A1(\cpuregs[9][15] ),
    .S(_19649_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _22801_ (.A0(_19625_),
    .A1(\cpuregs[9][14] ),
    .S(_19649_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _22802_ (.A(_19646_),
    .X(_19650_));
 sky130_fd_sc_hd__mux2_1 _22803_ (.A0(_19626_),
    .A1(\cpuregs[9][13] ),
    .S(_19650_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _22804_ (.A0(_19628_),
    .A1(\cpuregs[9][12] ),
    .S(_19650_),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _22805_ (.A0(_19629_),
    .A1(\cpuregs[9][11] ),
    .S(_19650_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _22806_ (.A0(_19630_),
    .A1(\cpuregs[9][10] ),
    .S(_19650_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _22807_ (.A0(_19631_),
    .A1(\cpuregs[9][9] ),
    .S(_19650_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _22808_ (.A0(_19632_),
    .A1(\cpuregs[9][8] ),
    .S(_19650_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_4 _22809_ (.A(_19645_),
    .X(_19651_));
 sky130_fd_sc_hd__mux2_1 _22810_ (.A0(_19633_),
    .A1(\cpuregs[9][7] ),
    .S(_19651_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _22811_ (.A0(_19635_),
    .A1(\cpuregs[9][6] ),
    .S(_19651_),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_1 _22812_ (.A0(_19636_),
    .A1(\cpuregs[9][5] ),
    .S(_19651_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _22813_ (.A0(_19637_),
    .A1(\cpuregs[9][4] ),
    .S(_19651_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _22814_ (.A0(_19638_),
    .A1(\cpuregs[9][3] ),
    .S(_19651_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _22815_ (.A0(_19639_),
    .A1(\cpuregs[9][2] ),
    .S(_19651_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _22816_ (.A0(_19640_),
    .A1(\cpuregs[9][1] ),
    .S(_19646_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _22817_ (.A0(_19641_),
    .A1(\cpuregs[9][0] ),
    .S(_19646_),
    .X(_03664_));
 sky130_fd_sc_hd__nor2_4 _22818_ (.A(_18533_),
    .B(_18959_),
    .Y(_19652_));
 sky130_fd_sc_hd__clkbuf_4 _22819_ (.A(_19652_),
    .X(_19653_));
 sky130_fd_sc_hd__buf_4 _22820_ (.A(_19653_),
    .X(_19654_));
 sky130_fd_sc_hd__mux2_1 _22821_ (.A0(net362),
    .A1(_02467_),
    .S(_19654_),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_1 _22822_ (.A0(net361),
    .A1(_02466_),
    .S(_19654_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_4 _22823_ (.A(net359),
    .X(_19655_));
 sky130_fd_sc_hd__mux2_1 _22824_ (.A0(_19655_),
    .A1(_02464_),
    .S(_19654_),
    .X(_03661_));
 sky130_fd_sc_hd__mux2_1 _22825_ (.A0(net358),
    .A1(_02463_),
    .S(_19654_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_4 _22826_ (.A(net357),
    .X(_19656_));
 sky130_fd_sc_hd__mux2_1 _22827_ (.A0(_19656_),
    .A1(_02462_),
    .S(_19654_),
    .X(_03659_));
 sky130_fd_sc_hd__buf_4 _22828_ (.A(net356),
    .X(_19657_));
 sky130_fd_sc_hd__buf_2 _22829_ (.A(_19653_),
    .X(_19658_));
 sky130_fd_sc_hd__mux2_1 _22830_ (.A0(_19657_),
    .A1(_02461_),
    .S(_19658_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_4 _22831_ (.A(net355),
    .X(_19659_));
 sky130_fd_sc_hd__mux2_1 _22832_ (.A0(_19659_),
    .A1(_02460_),
    .S(_19658_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _22833_ (.A0(net354),
    .A1(_02459_),
    .S(_19658_),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _22834_ (.A0(net353),
    .A1(_02458_),
    .S(_19658_),
    .X(_03655_));
 sky130_fd_sc_hd__mux2_1 _22835_ (.A0(net352),
    .A1(_02457_),
    .S(_19658_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_4 _22836_ (.A(net351),
    .X(_19660_));
 sky130_fd_sc_hd__mux2_1 _22837_ (.A0(_19660_),
    .A1(_02456_),
    .S(_19658_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_4 _22838_ (.A(_19653_),
    .X(_19661_));
 sky130_fd_sc_hd__mux2_1 _22839_ (.A0(net350),
    .A1(_02455_),
    .S(_19661_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _22840_ (.A0(net348),
    .A1(_02453_),
    .S(_19661_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_4 _22841_ (.A(net347),
    .X(_19662_));
 sky130_fd_sc_hd__mux2_1 _22842_ (.A0(_19662_),
    .A1(_02452_),
    .S(_19661_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_4 _22843_ (.A(net346),
    .X(_19663_));
 sky130_fd_sc_hd__mux2_1 _22844_ (.A0(_19663_),
    .A1(_02451_),
    .S(_19661_),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_1 _22845_ (.A0(net345),
    .A1(_02450_),
    .S(_19661_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_4 _22846_ (.A(net344),
    .X(_19664_));
 sky130_fd_sc_hd__mux2_1 _22847_ (.A0(_19664_),
    .A1(_02449_),
    .S(_19661_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_4 _22848_ (.A(_19652_),
    .X(_19665_));
 sky130_fd_sc_hd__mux2_1 _22849_ (.A0(net343),
    .A1(_02448_),
    .S(_19665_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_4 _22850_ (.A(net342),
    .X(_19666_));
 sky130_fd_sc_hd__mux2_1 _22851_ (.A0(_19666_),
    .A1(_02447_),
    .S(_19665_),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_1 _22852_ (.A0(net341),
    .A1(_02446_),
    .S(_19665_),
    .X(_03644_));
 sky130_fd_sc_hd__clkbuf_4 _22853_ (.A(net340),
    .X(_19667_));
 sky130_fd_sc_hd__mux2_1 _22854_ (.A0(_19667_),
    .A1(_02445_),
    .S(_19665_),
    .X(_03643_));
 sky130_fd_sc_hd__mux2_1 _22855_ (.A0(net339),
    .A1(_02444_),
    .S(_19665_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_2 _22856_ (.A(net369),
    .X(_19668_));
 sky130_fd_sc_hd__mux2_1 _22857_ (.A0(_19668_),
    .A1(_02474_),
    .S(_19665_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_2 _22858_ (.A(_19652_),
    .X(_19669_));
 sky130_fd_sc_hd__mux2_1 _22859_ (.A0(net368),
    .A1(_02473_),
    .S(_19669_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_8 _22860_ (.A(net229),
    .X(_19670_));
 sky130_fd_sc_hd__mux2_1 _22861_ (.A0(_19670_),
    .A1(_02472_),
    .S(_19669_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_6 _22862_ (.A(net228),
    .X(_19671_));
 sky130_fd_sc_hd__mux2_1 _22863_ (.A0(_19671_),
    .A1(_02471_),
    .S(_19669_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_6 _22864_ (.A(net227),
    .X(_19672_));
 sky130_fd_sc_hd__mux2_1 _22865_ (.A0(_19672_),
    .A1(_02470_),
    .S(_19669_),
    .X(_03637_));
 sky130_fd_sc_hd__buf_8 _22866_ (.A(net226),
    .X(_19673_));
 sky130_fd_sc_hd__mux2_1 _22867_ (.A0(_19673_),
    .A1(_02469_),
    .S(_19669_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_6 _22868_ (.A(net225),
    .X(_19674_));
 sky130_fd_sc_hd__mux2_1 _22869_ (.A0(_19674_),
    .A1(_02468_),
    .S(_19669_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_6 _22870_ (.A(net222),
    .X(_19675_));
 sky130_fd_sc_hd__mux2_1 _22871_ (.A0(_19675_),
    .A1(_02465_),
    .S(_19653_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_6 _22872_ (.A(net211),
    .X(_19676_));
 sky130_fd_sc_hd__mux2_1 _22873_ (.A0(_19676_),
    .A1(_02454_),
    .S(_19653_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_4 _22874_ (.A(net200),
    .X(_19677_));
 sky130_fd_sc_hd__mux2_1 _22875_ (.A0(_19677_),
    .A1(_02443_),
    .S(_19653_),
    .X(_03632_));
 sky130_fd_sc_hd__or3b_1 _22876_ (.A(_19592_),
    .B(_19599_),
    .C_N(_19603_),
    .X(_19678_));
 sky130_fd_sc_hd__buf_6 _22877_ (.A(_19678_),
    .X(_19679_));
 sky130_fd_sc_hd__clkbuf_4 _22878_ (.A(_19679_),
    .X(_19680_));
 sky130_fd_sc_hd__mux2_1 _22879_ (.A0(_19589_),
    .A1(\cpuregs[4][31] ),
    .S(_19680_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _22880_ (.A0(_19607_),
    .A1(\cpuregs[4][30] ),
    .S(_19680_),
    .X(_03630_));
 sky130_fd_sc_hd__mux2_1 _22881_ (.A0(_19608_),
    .A1(\cpuregs[4][29] ),
    .S(_19680_),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_1 _22882_ (.A0(_19609_),
    .A1(\cpuregs[4][28] ),
    .S(_19680_),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _22883_ (.A0(_19610_),
    .A1(\cpuregs[4][27] ),
    .S(_19680_),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_1 _22884_ (.A0(_19611_),
    .A1(\cpuregs[4][26] ),
    .S(_19680_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_4 _22885_ (.A(_19679_),
    .X(_19681_));
 sky130_fd_sc_hd__mux2_1 _22886_ (.A0(_19612_),
    .A1(\cpuregs[4][25] ),
    .S(_19681_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _22887_ (.A0(_19614_),
    .A1(\cpuregs[4][24] ),
    .S(_19681_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _22888_ (.A0(_19615_),
    .A1(\cpuregs[4][23] ),
    .S(_19681_),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_1 _22889_ (.A0(_19616_),
    .A1(\cpuregs[4][22] ),
    .S(_19681_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _22890_ (.A0(_19617_),
    .A1(\cpuregs[4][21] ),
    .S(_19681_),
    .X(_03621_));
 sky130_fd_sc_hd__mux2_1 _22891_ (.A0(_19618_),
    .A1(\cpuregs[4][20] ),
    .S(_19681_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_2 _22892_ (.A(_19679_),
    .X(_19682_));
 sky130_fd_sc_hd__mux2_1 _22893_ (.A0(_19619_),
    .A1(\cpuregs[4][19] ),
    .S(_19682_),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_1 _22894_ (.A0(_19621_),
    .A1(\cpuregs[4][18] ),
    .S(_19682_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _22895_ (.A0(_19622_),
    .A1(\cpuregs[4][17] ),
    .S(_19682_),
    .X(_03617_));
 sky130_fd_sc_hd__mux2_1 _22896_ (.A0(_19623_),
    .A1(\cpuregs[4][16] ),
    .S(_19682_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _22897_ (.A0(_19624_),
    .A1(\cpuregs[4][15] ),
    .S(_19682_),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_1 _22898_ (.A0(_19625_),
    .A1(\cpuregs[4][14] ),
    .S(_19682_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_4 _22899_ (.A(_19679_),
    .X(_19683_));
 sky130_fd_sc_hd__mux2_1 _22900_ (.A0(_19626_),
    .A1(\cpuregs[4][13] ),
    .S(_19683_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _22901_ (.A0(_19628_),
    .A1(\cpuregs[4][12] ),
    .S(_19683_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _22902_ (.A0(_19629_),
    .A1(\cpuregs[4][11] ),
    .S(_19683_),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_1 _22903_ (.A0(_19630_),
    .A1(\cpuregs[4][10] ),
    .S(_19683_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _22904_ (.A0(_19631_),
    .A1(\cpuregs[4][9] ),
    .S(_19683_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _22905_ (.A0(_19632_),
    .A1(\cpuregs[4][8] ),
    .S(_19683_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_4 _22906_ (.A(_19678_),
    .X(_19684_));
 sky130_fd_sc_hd__mux2_1 _22907_ (.A0(_19633_),
    .A1(\cpuregs[4][7] ),
    .S(_19684_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _22908_ (.A0(_19635_),
    .A1(\cpuregs[4][6] ),
    .S(_19684_),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _22909_ (.A0(_19636_),
    .A1(\cpuregs[4][5] ),
    .S(_19684_),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_1 _22910_ (.A0(_19637_),
    .A1(\cpuregs[4][4] ),
    .S(_19684_),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _22911_ (.A0(_19638_),
    .A1(\cpuregs[4][3] ),
    .S(_19684_),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _22912_ (.A0(_19639_),
    .A1(\cpuregs[4][2] ),
    .S(_19684_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _22913_ (.A0(_19640_),
    .A1(\cpuregs[4][1] ),
    .S(_19679_),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _22914_ (.A0(_19641_),
    .A1(\cpuregs[4][0] ),
    .S(_19679_),
    .X(_03600_));
 sky130_fd_sc_hd__nor2_4 _22915_ (.A(_19591_),
    .B(_19600_),
    .Y(_19685_));
 sky130_vsdinv _22916_ (.A(\latched_rd[2] ),
    .Y(_19686_));
 sky130_fd_sc_hd__and3_1 _22917_ (.A(_19686_),
    .B(_19594_),
    .C(\latched_rd[4] ),
    .X(_19687_));
 sky130_fd_sc_hd__nand2_1 _22918_ (.A(_19685_),
    .B(_19687_),
    .Y(_19688_));
 sky130_fd_sc_hd__buf_4 _22919_ (.A(_19688_),
    .X(_19689_));
 sky130_fd_sc_hd__clkbuf_4 _22920_ (.A(_19689_),
    .X(_19690_));
 sky130_fd_sc_hd__mux2_1 _22921_ (.A0(_19589_),
    .A1(\cpuregs[19][31] ),
    .S(_19690_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _22922_ (.A0(_19607_),
    .A1(\cpuregs[19][30] ),
    .S(_19690_),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_1 _22923_ (.A0(_19608_),
    .A1(\cpuregs[19][29] ),
    .S(_19690_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _22924_ (.A0(_19609_),
    .A1(\cpuregs[19][28] ),
    .S(_19690_),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_1 _22925_ (.A0(_19610_),
    .A1(\cpuregs[19][27] ),
    .S(_19690_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_1 _22926_ (.A0(_19611_),
    .A1(\cpuregs[19][26] ),
    .S(_19690_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_4 _22927_ (.A(_19689_),
    .X(_19691_));
 sky130_fd_sc_hd__mux2_1 _22928_ (.A0(_19612_),
    .A1(\cpuregs[19][25] ),
    .S(_19691_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _22929_ (.A0(_19614_),
    .A1(\cpuregs[19][24] ),
    .S(_19691_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _22930_ (.A0(_19615_),
    .A1(\cpuregs[19][23] ),
    .S(_19691_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _22931_ (.A0(_19616_),
    .A1(\cpuregs[19][22] ),
    .S(_19691_),
    .X(_03590_));
 sky130_fd_sc_hd__mux2_1 _22932_ (.A0(_19617_),
    .A1(\cpuregs[19][21] ),
    .S(_19691_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _22933_ (.A0(_19618_),
    .A1(\cpuregs[19][20] ),
    .S(_19691_),
    .X(_03588_));
 sky130_fd_sc_hd__buf_2 _22934_ (.A(_19689_),
    .X(_19692_));
 sky130_fd_sc_hd__mux2_1 _22935_ (.A0(_19619_),
    .A1(\cpuregs[19][19] ),
    .S(_19692_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _22936_ (.A0(_19621_),
    .A1(\cpuregs[19][18] ),
    .S(_19692_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_1 _22937_ (.A0(_19622_),
    .A1(\cpuregs[19][17] ),
    .S(_19692_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _22938_ (.A0(_19623_),
    .A1(\cpuregs[19][16] ),
    .S(_19692_),
    .X(_03584_));
 sky130_fd_sc_hd__mux2_1 _22939_ (.A0(_19624_),
    .A1(\cpuregs[19][15] ),
    .S(_19692_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _22940_ (.A0(_19625_),
    .A1(\cpuregs[19][14] ),
    .S(_19692_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_4 _22941_ (.A(_19689_),
    .X(_19693_));
 sky130_fd_sc_hd__mux2_1 _22942_ (.A0(_19626_),
    .A1(\cpuregs[19][13] ),
    .S(_19693_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _22943_ (.A0(_19628_),
    .A1(\cpuregs[19][12] ),
    .S(_19693_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_1 _22944_ (.A0(_19629_),
    .A1(\cpuregs[19][11] ),
    .S(_19693_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_1 _22945_ (.A0(_19630_),
    .A1(\cpuregs[19][10] ),
    .S(_19693_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_1 _22946_ (.A0(_19631_),
    .A1(\cpuregs[19][9] ),
    .S(_19693_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _22947_ (.A0(_19632_),
    .A1(\cpuregs[19][8] ),
    .S(_19693_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_4 _22948_ (.A(_19688_),
    .X(_19694_));
 sky130_fd_sc_hd__mux2_1 _22949_ (.A0(_19633_),
    .A1(\cpuregs[19][7] ),
    .S(_19694_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _22950_ (.A0(_19635_),
    .A1(\cpuregs[19][6] ),
    .S(_19694_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _22951_ (.A0(_19636_),
    .A1(\cpuregs[19][5] ),
    .S(_19694_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _22952_ (.A0(_19637_),
    .A1(\cpuregs[19][4] ),
    .S(_19694_),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_1 _22953_ (.A0(_19638_),
    .A1(\cpuregs[19][3] ),
    .S(_19694_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _22954_ (.A0(_19639_),
    .A1(\cpuregs[19][2] ),
    .S(_19694_),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_1 _22955_ (.A0(_19640_),
    .A1(\cpuregs[19][1] ),
    .S(_19689_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _22956_ (.A0(_19641_),
    .A1(\cpuregs[19][0] ),
    .S(_19689_),
    .X(_03568_));
 sky130_fd_sc_hd__nand2_1 _22957_ (.A(_18855_),
    .B(mem_do_wdata),
    .Y(_19695_));
 sky130_fd_sc_hd__or2_4 _22958_ (.A(net408),
    .B(_19695_),
    .X(_19696_));
 sky130_fd_sc_hd__clkbuf_2 _22959_ (.A(_19696_),
    .X(_19697_));
 sky130_fd_sc_hd__buf_4 _22960_ (.A(_19697_),
    .X(_19698_));
 sky130_fd_sc_hd__mux2_1 _22961_ (.A0(net224),
    .A1(net262),
    .S(net424),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_1 _22962_ (.A0(net223),
    .A1(net261),
    .S(net424),
    .X(_03566_));
 sky130_fd_sc_hd__mux2_1 _22963_ (.A0(net221),
    .A1(net259),
    .S(net424),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_1 _22964_ (.A0(net220),
    .A1(net258),
    .S(net424),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_1 _22965_ (.A0(net219),
    .A1(net257),
    .S(_19698_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _22966_ (.A0(net218),
    .A1(net256),
    .S(net424),
    .X(_03562_));
 sky130_fd_sc_hd__buf_6 _22967_ (.A(_19697_),
    .X(_19699_));
 sky130_fd_sc_hd__mux2_1 _22968_ (.A0(net217),
    .A1(net255),
    .S(_19699_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _22969_ (.A0(net216),
    .A1(net254),
    .S(_19699_),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _22970_ (.A0(net215),
    .A1(net253),
    .S(_19699_),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_1 _22971_ (.A0(net214),
    .A1(net252),
    .S(_19699_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _22972_ (.A0(net213),
    .A1(net251),
    .S(_19699_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _22973_ (.A0(net212),
    .A1(net250),
    .S(_19699_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_4 _22974_ (.A(_19697_),
    .X(_19700_));
 sky130_fd_sc_hd__mux2_1 _22975_ (.A0(net210),
    .A1(net248),
    .S(net422),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_1 _22976_ (.A0(net209),
    .A1(net247),
    .S(net422),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_1 _22977_ (.A0(net208),
    .A1(net246),
    .S(net423),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_1 _22978_ (.A0(net207),
    .A1(net245),
    .S(_19700_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _22979_ (.A0(net206),
    .A1(net244),
    .S(net422),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_1 _22980_ (.A0(net205),
    .A1(net243),
    .S(net423),
    .X(_03550_));
 sky130_fd_sc_hd__buf_4 _22981_ (.A(_19697_),
    .X(_19701_));
 sky130_fd_sc_hd__mux2_1 _22982_ (.A0(net204),
    .A1(net242),
    .S(net421),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _22983_ (.A0(net203),
    .A1(net241),
    .S(_19701_),
    .X(_03548_));
 sky130_fd_sc_hd__mux2_1 _22984_ (.A0(net202),
    .A1(net240),
    .S(_19701_),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_1 _22985_ (.A0(net201),
    .A1(net239),
    .S(_19701_),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _22986_ (.A0(net231),
    .A1(net269),
    .S(net421),
    .X(_03545_));
 sky130_fd_sc_hd__mux2_1 _22987_ (.A0(net230),
    .A1(net268),
    .S(net421),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_2 _22988_ (.A(_19696_),
    .X(_19702_));
 sky130_fd_sc_hd__mux2_1 _22989_ (.A0(_19670_),
    .A1(net267),
    .S(net426),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _22990_ (.A0(_19671_),
    .A1(net266),
    .S(net426),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_1 _22991_ (.A0(_19672_),
    .A1(net265),
    .S(_19702_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _22992_ (.A0(_19673_),
    .A1(net264),
    .S(net426),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_1 _22993_ (.A0(_19674_),
    .A1(net263),
    .S(_19702_),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _22994_ (.A0(_19675_),
    .A1(net260),
    .S(net426),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_1 _22995_ (.A0(_19676_),
    .A1(net249),
    .S(_19697_),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_1 _22996_ (.A0(_19677_),
    .A1(net238),
    .S(_19697_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_1 _22997_ (.A(_19685_),
    .B(_19603_),
    .Y(_19703_));
 sky130_fd_sc_hd__buf_6 _22998_ (.A(_19703_),
    .X(_19704_));
 sky130_fd_sc_hd__clkbuf_4 _22999_ (.A(_19704_),
    .X(_19705_));
 sky130_fd_sc_hd__mux2_1 _23000_ (.A0(_19589_),
    .A1(\cpuregs[7][31] ),
    .S(_19705_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_1 _23001_ (.A0(_19607_),
    .A1(\cpuregs[7][30] ),
    .S(_19705_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _23002_ (.A0(_19608_),
    .A1(\cpuregs[7][29] ),
    .S(_19705_),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_1 _23003_ (.A0(_19609_),
    .A1(\cpuregs[7][28] ),
    .S(_19705_),
    .X(_03532_));
 sky130_fd_sc_hd__mux2_1 _23004_ (.A0(_19610_),
    .A1(\cpuregs[7][27] ),
    .S(_19705_),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_1 _23005_ (.A0(_19611_),
    .A1(\cpuregs[7][26] ),
    .S(_19705_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_4 _23006_ (.A(_19704_),
    .X(_19706_));
 sky130_fd_sc_hd__mux2_1 _23007_ (.A0(_19612_),
    .A1(\cpuregs[7][25] ),
    .S(_19706_),
    .X(_03529_));
 sky130_fd_sc_hd__mux2_1 _23008_ (.A0(_19614_),
    .A1(\cpuregs[7][24] ),
    .S(_19706_),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_1 _23009_ (.A0(_19615_),
    .A1(\cpuregs[7][23] ),
    .S(_19706_),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_1 _23010_ (.A0(_19616_),
    .A1(\cpuregs[7][22] ),
    .S(_19706_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_1 _23011_ (.A0(_19617_),
    .A1(\cpuregs[7][21] ),
    .S(_19706_),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_1 _23012_ (.A0(_19618_),
    .A1(\cpuregs[7][20] ),
    .S(_19706_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_4 _23013_ (.A(_19704_),
    .X(_19707_));
 sky130_fd_sc_hd__mux2_1 _23014_ (.A0(_19619_),
    .A1(\cpuregs[7][19] ),
    .S(_19707_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _23015_ (.A0(_19621_),
    .A1(\cpuregs[7][18] ),
    .S(_19707_),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_1 _23016_ (.A0(_19622_),
    .A1(\cpuregs[7][17] ),
    .S(_19707_),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_1 _23017_ (.A0(_19623_),
    .A1(\cpuregs[7][16] ),
    .S(_19707_),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _23018_ (.A0(_19624_),
    .A1(\cpuregs[7][15] ),
    .S(_19707_),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_1 _23019_ (.A0(_19625_),
    .A1(\cpuregs[7][14] ),
    .S(_19707_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_4 _23020_ (.A(_19704_),
    .X(_19708_));
 sky130_fd_sc_hd__mux2_1 _23021_ (.A0(_19626_),
    .A1(\cpuregs[7][13] ),
    .S(_19708_),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_1 _23022_ (.A0(_19628_),
    .A1(\cpuregs[7][12] ),
    .S(_19708_),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_1 _23023_ (.A0(_19629_),
    .A1(\cpuregs[7][11] ),
    .S(_19708_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_1 _23024_ (.A0(_19630_),
    .A1(\cpuregs[7][10] ),
    .S(_19708_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _23025_ (.A0(_19631_),
    .A1(\cpuregs[7][9] ),
    .S(_19708_),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_1 _23026_ (.A0(_19632_),
    .A1(\cpuregs[7][8] ),
    .S(_19708_),
    .X(_03512_));
 sky130_fd_sc_hd__clkbuf_4 _23027_ (.A(_19703_),
    .X(_19709_));
 sky130_fd_sc_hd__mux2_1 _23028_ (.A0(_19633_),
    .A1(\cpuregs[7][7] ),
    .S(_19709_),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _23029_ (.A0(_19635_),
    .A1(\cpuregs[7][6] ),
    .S(_19709_),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_1 _23030_ (.A0(_19636_),
    .A1(\cpuregs[7][5] ),
    .S(_19709_),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _23031_ (.A0(_19637_),
    .A1(\cpuregs[7][4] ),
    .S(_19709_),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_1 _23032_ (.A0(_19638_),
    .A1(\cpuregs[7][3] ),
    .S(_19709_),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_1 _23033_ (.A0(_19639_),
    .A1(\cpuregs[7][2] ),
    .S(_19709_),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_1 _23034_ (.A0(_19640_),
    .A1(\cpuregs[7][1] ),
    .S(_19704_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _23035_ (.A0(_19641_),
    .A1(\cpuregs[7][0] ),
    .S(_19704_),
    .X(_03504_));
 sky130_fd_sc_hd__nand2_1 _23036_ (.A(_18768_),
    .B(_18700_),
    .Y(_19710_));
 sky130_fd_sc_hd__o2111a_1 _23037_ (.A1(instr_setq),
    .A2(_19316_),
    .B1(_18547_),
    .C1(_18553_),
    .D1(_19710_),
    .X(_19711_));
 sky130_fd_sc_hd__mux2_1 _23038_ (.A0(\latched_rd[4] ),
    .A1(_21104_),
    .S(_19711_),
    .X(_03503_));
 sky130_fd_sc_hd__and3_1 _23039_ (.A(_19602_),
    .B(\latched_rd[2] ),
    .C(\latched_rd[3] ),
    .X(_19712_));
 sky130_fd_sc_hd__nand2_1 _23040_ (.A(_19685_),
    .B(_19712_),
    .Y(_19713_));
 sky130_fd_sc_hd__buf_6 _23041_ (.A(_19713_),
    .X(_19714_));
 sky130_fd_sc_hd__clkbuf_4 _23042_ (.A(_19714_),
    .X(_19715_));
 sky130_fd_sc_hd__mux2_1 _23043_ (.A0(_19589_),
    .A1(\cpuregs[15][31] ),
    .S(_19715_),
    .X(_03502_));
 sky130_fd_sc_hd__mux2_1 _23044_ (.A0(_19607_),
    .A1(\cpuregs[15][30] ),
    .S(_19715_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _23045_ (.A0(_19608_),
    .A1(\cpuregs[15][29] ),
    .S(_19715_),
    .X(_03500_));
 sky130_fd_sc_hd__mux2_1 _23046_ (.A0(_19609_),
    .A1(\cpuregs[15][28] ),
    .S(_19715_),
    .X(_03499_));
 sky130_fd_sc_hd__mux2_1 _23047_ (.A0(_19610_),
    .A1(\cpuregs[15][27] ),
    .S(_19715_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_1 _23048_ (.A0(_19611_),
    .A1(\cpuregs[15][26] ),
    .S(_19715_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_4 _23049_ (.A(_19714_),
    .X(_19716_));
 sky130_fd_sc_hd__mux2_1 _23050_ (.A0(_19612_),
    .A1(\cpuregs[15][25] ),
    .S(_19716_),
    .X(_03496_));
 sky130_fd_sc_hd__mux2_1 _23051_ (.A0(_19614_),
    .A1(\cpuregs[15][24] ),
    .S(_19716_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _23052_ (.A0(_19615_),
    .A1(\cpuregs[15][23] ),
    .S(_19716_),
    .X(_03494_));
 sky130_fd_sc_hd__mux2_1 _23053_ (.A0(_19616_),
    .A1(\cpuregs[15][22] ),
    .S(_19716_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_1 _23054_ (.A0(_19617_),
    .A1(\cpuregs[15][21] ),
    .S(_19716_),
    .X(_03492_));
 sky130_fd_sc_hd__mux2_1 _23055_ (.A0(_19618_),
    .A1(\cpuregs[15][20] ),
    .S(_19716_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_4 _23056_ (.A(_19714_),
    .X(_19717_));
 sky130_fd_sc_hd__mux2_1 _23057_ (.A0(_19619_),
    .A1(\cpuregs[15][19] ),
    .S(_19717_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _23058_ (.A0(_19621_),
    .A1(\cpuregs[15][18] ),
    .S(_19717_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _23059_ (.A0(_19622_),
    .A1(\cpuregs[15][17] ),
    .S(_19717_),
    .X(_03488_));
 sky130_fd_sc_hd__mux2_1 _23060_ (.A0(_19623_),
    .A1(\cpuregs[15][16] ),
    .S(_19717_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _23061_ (.A0(_19624_),
    .A1(\cpuregs[15][15] ),
    .S(_19717_),
    .X(_03486_));
 sky130_fd_sc_hd__mux2_1 _23062_ (.A0(_19625_),
    .A1(\cpuregs[15][14] ),
    .S(_19717_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_4 _23063_ (.A(_19714_),
    .X(_19718_));
 sky130_fd_sc_hd__mux2_1 _23064_ (.A0(_19626_),
    .A1(\cpuregs[15][13] ),
    .S(_19718_),
    .X(_03484_));
 sky130_fd_sc_hd__mux2_1 _23065_ (.A0(_19628_),
    .A1(\cpuregs[15][12] ),
    .S(_19718_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _23066_ (.A0(_19629_),
    .A1(\cpuregs[15][11] ),
    .S(_19718_),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_1 _23067_ (.A0(_19630_),
    .A1(\cpuregs[15][10] ),
    .S(_19718_),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _23068_ (.A0(_19631_),
    .A1(\cpuregs[15][9] ),
    .S(_19718_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _23069_ (.A0(_19632_),
    .A1(\cpuregs[15][8] ),
    .S(_19718_),
    .X(_03479_));
 sky130_fd_sc_hd__buf_2 _23070_ (.A(_19713_),
    .X(_19719_));
 sky130_fd_sc_hd__mux2_1 _23071_ (.A0(_19633_),
    .A1(\cpuregs[15][7] ),
    .S(_19719_),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_1 _23072_ (.A0(_19635_),
    .A1(\cpuregs[15][6] ),
    .S(_19719_),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_1 _23073_ (.A0(_19636_),
    .A1(\cpuregs[15][5] ),
    .S(_19719_),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_1 _23074_ (.A0(_19637_),
    .A1(\cpuregs[15][4] ),
    .S(_19719_),
    .X(_03475_));
 sky130_fd_sc_hd__mux2_1 _23075_ (.A0(_19638_),
    .A1(\cpuregs[15][3] ),
    .S(_19719_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _23076_ (.A0(_19639_),
    .A1(\cpuregs[15][2] ),
    .S(_19719_),
    .X(_03473_));
 sky130_fd_sc_hd__mux2_1 _23077_ (.A0(_19640_),
    .A1(\cpuregs[15][1] ),
    .S(_19714_),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_1 _23078_ (.A0(_19641_),
    .A1(\cpuregs[15][0] ),
    .S(_19714_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_2 _23079_ (.A(\cpuregs_wrdata[31] ),
    .X(_19720_));
 sky130_fd_sc_hd__nand2_1 _23080_ (.A(_19685_),
    .B(_19644_),
    .Y(_19721_));
 sky130_fd_sc_hd__buf_6 _23081_ (.A(_19721_),
    .X(_19722_));
 sky130_fd_sc_hd__buf_4 _23082_ (.A(_19722_),
    .X(_19723_));
 sky130_fd_sc_hd__mux2_1 _23083_ (.A0(_19720_),
    .A1(\cpuregs[11][31] ),
    .S(_19723_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_2 _23084_ (.A(\cpuregs_wrdata[30] ),
    .X(_19724_));
 sky130_fd_sc_hd__mux2_1 _23085_ (.A0(_19724_),
    .A1(\cpuregs[11][30] ),
    .S(_19723_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_2 _23086_ (.A(\cpuregs_wrdata[29] ),
    .X(_19725_));
 sky130_fd_sc_hd__mux2_1 _23087_ (.A0(_19725_),
    .A1(\cpuregs[11][29] ),
    .S(_19723_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_2 _23088_ (.A(\cpuregs_wrdata[28] ),
    .X(_19726_));
 sky130_fd_sc_hd__mux2_1 _23089_ (.A0(_19726_),
    .A1(\cpuregs[11][28] ),
    .S(_19723_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_2 _23090_ (.A(\cpuregs_wrdata[27] ),
    .X(_19727_));
 sky130_fd_sc_hd__mux2_1 _23091_ (.A0(_19727_),
    .A1(\cpuregs[11][27] ),
    .S(_19723_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_2 _23092_ (.A(\cpuregs_wrdata[26] ),
    .X(_19728_));
 sky130_fd_sc_hd__mux2_1 _23093_ (.A0(_19728_),
    .A1(\cpuregs[11][26] ),
    .S(_19723_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_2 _23094_ (.A(\cpuregs_wrdata[25] ),
    .X(_19729_));
 sky130_fd_sc_hd__clkbuf_4 _23095_ (.A(_19722_),
    .X(_19730_));
 sky130_fd_sc_hd__mux2_1 _23096_ (.A0(_19729_),
    .A1(\cpuregs[11][25] ),
    .S(_19730_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_2 _23097_ (.A(\cpuregs_wrdata[24] ),
    .X(_19731_));
 sky130_fd_sc_hd__mux2_1 _23098_ (.A0(_19731_),
    .A1(\cpuregs[11][24] ),
    .S(_19730_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_2 _23099_ (.A(\cpuregs_wrdata[23] ),
    .X(_19732_));
 sky130_fd_sc_hd__mux2_1 _23100_ (.A0(_19732_),
    .A1(\cpuregs[11][23] ),
    .S(_19730_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_2 _23101_ (.A(\cpuregs_wrdata[22] ),
    .X(_19733_));
 sky130_fd_sc_hd__mux2_1 _23102_ (.A0(_19733_),
    .A1(\cpuregs[11][22] ),
    .S(_19730_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_2 _23103_ (.A(\cpuregs_wrdata[21] ),
    .X(_19734_));
 sky130_fd_sc_hd__mux2_1 _23104_ (.A0(_19734_),
    .A1(\cpuregs[11][21] ),
    .S(_19730_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_2 _23105_ (.A(\cpuregs_wrdata[20] ),
    .X(_19735_));
 sky130_fd_sc_hd__mux2_1 _23106_ (.A0(_19735_),
    .A1(\cpuregs[11][20] ),
    .S(_19730_),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_2 _23107_ (.A(\cpuregs_wrdata[19] ),
    .X(_19736_));
 sky130_fd_sc_hd__clkbuf_4 _23108_ (.A(_19722_),
    .X(_19737_));
 sky130_fd_sc_hd__mux2_1 _23109_ (.A0(_19736_),
    .A1(\cpuregs[11][19] ),
    .S(_19737_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_2 _23110_ (.A(\cpuregs_wrdata[18] ),
    .X(_19738_));
 sky130_fd_sc_hd__mux2_1 _23111_ (.A0(_19738_),
    .A1(\cpuregs[11][18] ),
    .S(_19737_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_2 _23112_ (.A(\cpuregs_wrdata[17] ),
    .X(_19739_));
 sky130_fd_sc_hd__mux2_1 _23113_ (.A0(_19739_),
    .A1(\cpuregs[11][17] ),
    .S(_19737_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_2 _23114_ (.A(\cpuregs_wrdata[16] ),
    .X(_19740_));
 sky130_fd_sc_hd__mux2_1 _23115_ (.A0(_19740_),
    .A1(\cpuregs[11][16] ),
    .S(_19737_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_2 _23116_ (.A(\cpuregs_wrdata[15] ),
    .X(_19741_));
 sky130_fd_sc_hd__mux2_1 _23117_ (.A0(_19741_),
    .A1(\cpuregs[11][15] ),
    .S(_19737_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_2 _23118_ (.A(\cpuregs_wrdata[14] ),
    .X(_19742_));
 sky130_fd_sc_hd__mux2_1 _23119_ (.A0(_19742_),
    .A1(\cpuregs[11][14] ),
    .S(_19737_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_2 _23120_ (.A(\cpuregs_wrdata[13] ),
    .X(_19743_));
 sky130_fd_sc_hd__clkbuf_4 _23121_ (.A(_19722_),
    .X(_19744_));
 sky130_fd_sc_hd__mux2_1 _23122_ (.A0(_19743_),
    .A1(\cpuregs[11][13] ),
    .S(_19744_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_2 _23123_ (.A(\cpuregs_wrdata[12] ),
    .X(_19745_));
 sky130_fd_sc_hd__mux2_1 _23124_ (.A0(_19745_),
    .A1(\cpuregs[11][12] ),
    .S(_19744_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_2 _23125_ (.A(\cpuregs_wrdata[11] ),
    .X(_19746_));
 sky130_fd_sc_hd__mux2_1 _23126_ (.A0(_19746_),
    .A1(\cpuregs[11][11] ),
    .S(_19744_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_2 _23127_ (.A(\cpuregs_wrdata[10] ),
    .X(_19747_));
 sky130_fd_sc_hd__mux2_1 _23128_ (.A0(_19747_),
    .A1(\cpuregs[11][10] ),
    .S(_19744_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_2 _23129_ (.A(\cpuregs_wrdata[9] ),
    .X(_19748_));
 sky130_fd_sc_hd__mux2_1 _23130_ (.A0(_19748_),
    .A1(\cpuregs[11][9] ),
    .S(_19744_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_2 _23131_ (.A(\cpuregs_wrdata[8] ),
    .X(_19749_));
 sky130_fd_sc_hd__mux2_1 _23132_ (.A0(_19749_),
    .A1(\cpuregs[11][8] ),
    .S(_19744_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_2 _23133_ (.A(\cpuregs_wrdata[7] ),
    .X(_19750_));
 sky130_fd_sc_hd__clkbuf_4 _23134_ (.A(_19721_),
    .X(_19751_));
 sky130_fd_sc_hd__mux2_1 _23135_ (.A0(_19750_),
    .A1(\cpuregs[11][7] ),
    .S(_19751_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_2 _23136_ (.A(\cpuregs_wrdata[6] ),
    .X(_19752_));
 sky130_fd_sc_hd__mux2_1 _23137_ (.A0(_19752_),
    .A1(\cpuregs[11][6] ),
    .S(_19751_),
    .X(_03445_));
 sky130_fd_sc_hd__buf_2 _23138_ (.A(\cpuregs_wrdata[5] ),
    .X(_19753_));
 sky130_fd_sc_hd__mux2_1 _23139_ (.A0(_19753_),
    .A1(\cpuregs[11][5] ),
    .S(_19751_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_2 _23140_ (.A(\cpuregs_wrdata[4] ),
    .X(_19754_));
 sky130_fd_sc_hd__mux2_1 _23141_ (.A0(_19754_),
    .A1(\cpuregs[11][4] ),
    .S(_19751_),
    .X(_03443_));
 sky130_fd_sc_hd__clkbuf_2 _23142_ (.A(\cpuregs_wrdata[3] ),
    .X(_19755_));
 sky130_fd_sc_hd__mux2_1 _23143_ (.A0(_19755_),
    .A1(\cpuregs[11][3] ),
    .S(_19751_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_2 _23144_ (.A(\cpuregs_wrdata[2] ),
    .X(_19756_));
 sky130_fd_sc_hd__mux2_1 _23145_ (.A0(_19756_),
    .A1(\cpuregs[11][2] ),
    .S(_19751_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_2 _23146_ (.A(\cpuregs_wrdata[1] ),
    .X(_19757_));
 sky130_fd_sc_hd__mux2_1 _23147_ (.A0(_19757_),
    .A1(\cpuregs[11][1] ),
    .S(_19722_),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_2 _23148_ (.A(\cpuregs_wrdata[0] ),
    .X(_19758_));
 sky130_fd_sc_hd__mux2_1 _23149_ (.A0(_19758_),
    .A1(\cpuregs[11][0] ),
    .S(_19722_),
    .X(_03439_));
 sky130_vsdinv _23150_ (.A(_19595_),
    .Y(_19759_));
 sky130_fd_sc_hd__nand2_1 _23151_ (.A(_19685_),
    .B(_19759_),
    .Y(_19760_));
 sky130_fd_sc_hd__buf_6 _23152_ (.A(_19760_),
    .X(_19761_));
 sky130_fd_sc_hd__buf_4 _23153_ (.A(_19761_),
    .X(_19762_));
 sky130_fd_sc_hd__mux2_1 _23154_ (.A0(_19720_),
    .A1(\cpuregs[3][31] ),
    .S(_19762_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_1 _23155_ (.A0(_19724_),
    .A1(\cpuregs[3][30] ),
    .S(_19762_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _23156_ (.A0(_19725_),
    .A1(\cpuregs[3][29] ),
    .S(_19762_),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_1 _23157_ (.A0(_19726_),
    .A1(\cpuregs[3][28] ),
    .S(_19762_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _23158_ (.A0(_19727_),
    .A1(\cpuregs[3][27] ),
    .S(_19762_),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_1 _23159_ (.A0(_19728_),
    .A1(\cpuregs[3][26] ),
    .S(_19762_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_4 _23160_ (.A(_19761_),
    .X(_19763_));
 sky130_fd_sc_hd__mux2_1 _23161_ (.A0(_19729_),
    .A1(\cpuregs[3][25] ),
    .S(_19763_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _23162_ (.A0(_19731_),
    .A1(\cpuregs[3][24] ),
    .S(_19763_),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_1 _23163_ (.A0(_19732_),
    .A1(\cpuregs[3][23] ),
    .S(_19763_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_1 _23164_ (.A0(_19733_),
    .A1(\cpuregs[3][22] ),
    .S(_19763_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _23165_ (.A0(_19734_),
    .A1(\cpuregs[3][21] ),
    .S(_19763_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _23166_ (.A0(_19735_),
    .A1(\cpuregs[3][20] ),
    .S(_19763_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_4 _23167_ (.A(_19761_),
    .X(_19764_));
 sky130_fd_sc_hd__mux2_1 _23168_ (.A0(_19736_),
    .A1(\cpuregs[3][19] ),
    .S(_19764_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _23169_ (.A0(_19738_),
    .A1(\cpuregs[3][18] ),
    .S(_19764_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _23170_ (.A0(_19739_),
    .A1(\cpuregs[3][17] ),
    .S(_19764_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_1 _23171_ (.A0(_19740_),
    .A1(\cpuregs[3][16] ),
    .S(_19764_),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _23172_ (.A0(_19741_),
    .A1(\cpuregs[3][15] ),
    .S(_19764_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _23173_ (.A0(_19742_),
    .A1(\cpuregs[3][14] ),
    .S(_19764_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_4 _23174_ (.A(_19761_),
    .X(_19765_));
 sky130_fd_sc_hd__mux2_1 _23175_ (.A0(_19743_),
    .A1(\cpuregs[3][13] ),
    .S(_19765_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _23176_ (.A0(_19745_),
    .A1(\cpuregs[3][12] ),
    .S(_19765_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _23177_ (.A0(_19746_),
    .A1(\cpuregs[3][11] ),
    .S(_19765_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_1 _23178_ (.A0(_19747_),
    .A1(\cpuregs[3][10] ),
    .S(_19765_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _23179_ (.A0(_19748_),
    .A1(\cpuregs[3][9] ),
    .S(_19765_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_1 _23180_ (.A0(_19749_),
    .A1(\cpuregs[3][8] ),
    .S(_19765_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_4 _23181_ (.A(_19760_),
    .X(_19766_));
 sky130_fd_sc_hd__mux2_1 _23182_ (.A0(_19750_),
    .A1(\cpuregs[3][7] ),
    .S(_19766_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _23183_ (.A0(_19752_),
    .A1(\cpuregs[3][6] ),
    .S(_19766_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _23184_ (.A0(_19753_),
    .A1(\cpuregs[3][5] ),
    .S(_19766_),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_1 _23185_ (.A0(_19754_),
    .A1(\cpuregs[3][4] ),
    .S(_19766_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _23186_ (.A0(_19755_),
    .A1(\cpuregs[3][3] ),
    .S(_19766_),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_1 _23187_ (.A0(_19756_),
    .A1(\cpuregs[3][2] ),
    .S(_19766_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_1 _23188_ (.A0(_19757_),
    .A1(\cpuregs[3][1] ),
    .S(_19761_),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_1 _23189_ (.A0(_19758_),
    .A1(\cpuregs[3][0] ),
    .S(_19761_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_2 _23190_ (.A(\cpuregs_wrdata[31] ),
    .X(_19767_));
 sky130_fd_sc_hd__and2_1 _23191_ (.A(_19642_),
    .B(_19759_),
    .X(_19768_));
 sky130_fd_sc_hd__buf_6 _23192_ (.A(_19768_),
    .X(_19769_));
 sky130_fd_sc_hd__buf_4 _23193_ (.A(_19769_),
    .X(_19770_));
 sky130_fd_sc_hd__mux2_1 _23194_ (.A0(\cpuregs[1][31] ),
    .A1(_19767_),
    .S(_19770_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_2 _23195_ (.A(\cpuregs_wrdata[30] ),
    .X(_19771_));
 sky130_fd_sc_hd__mux2_1 _23196_ (.A0(\cpuregs[1][30] ),
    .A1(_19771_),
    .S(_19770_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_2 _23197_ (.A(\cpuregs_wrdata[29] ),
    .X(_19772_));
 sky130_fd_sc_hd__mux2_1 _23198_ (.A0(\cpuregs[1][29] ),
    .A1(_19772_),
    .S(_19770_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_2 _23199_ (.A(\cpuregs_wrdata[28] ),
    .X(_19773_));
 sky130_fd_sc_hd__mux2_1 _23200_ (.A0(\cpuregs[1][28] ),
    .A1(_19773_),
    .S(_19770_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_2 _23201_ (.A(\cpuregs_wrdata[27] ),
    .X(_19774_));
 sky130_fd_sc_hd__mux2_1 _23202_ (.A0(\cpuregs[1][27] ),
    .A1(_19774_),
    .S(_19770_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_2 _23203_ (.A(\cpuregs_wrdata[26] ),
    .X(_19775_));
 sky130_fd_sc_hd__mux2_1 _23204_ (.A0(\cpuregs[1][26] ),
    .A1(_19775_),
    .S(_19770_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_2 _23205_ (.A(\cpuregs_wrdata[25] ),
    .X(_19776_));
 sky130_fd_sc_hd__buf_4 _23206_ (.A(_19769_),
    .X(_19777_));
 sky130_fd_sc_hd__mux2_1 _23207_ (.A0(\cpuregs[1][25] ),
    .A1(_19776_),
    .S(_19777_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_2 _23208_ (.A(\cpuregs_wrdata[24] ),
    .X(_19778_));
 sky130_fd_sc_hd__mux2_1 _23209_ (.A0(\cpuregs[1][24] ),
    .A1(_19778_),
    .S(_19777_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_2 _23210_ (.A(\cpuregs_wrdata[23] ),
    .X(_19779_));
 sky130_fd_sc_hd__mux2_1 _23211_ (.A0(\cpuregs[1][23] ),
    .A1(_19779_),
    .S(_19777_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_2 _23212_ (.A(\cpuregs_wrdata[22] ),
    .X(_19780_));
 sky130_fd_sc_hd__mux2_1 _23213_ (.A0(\cpuregs[1][22] ),
    .A1(_19780_),
    .S(_19777_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_2 _23214_ (.A(\cpuregs_wrdata[21] ),
    .X(_19781_));
 sky130_fd_sc_hd__mux2_1 _23215_ (.A0(\cpuregs[1][21] ),
    .A1(_19781_),
    .S(_19777_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_2 _23216_ (.A(\cpuregs_wrdata[20] ),
    .X(_19782_));
 sky130_fd_sc_hd__mux2_1 _23217_ (.A0(\cpuregs[1][20] ),
    .A1(_19782_),
    .S(_19777_),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_2 _23218_ (.A(\cpuregs_wrdata[19] ),
    .X(_19783_));
 sky130_fd_sc_hd__clkbuf_4 _23219_ (.A(_19769_),
    .X(_19784_));
 sky130_fd_sc_hd__mux2_1 _23220_ (.A0(\cpuregs[1][19] ),
    .A1(_19783_),
    .S(_19784_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_2 _23221_ (.A(\cpuregs_wrdata[18] ),
    .X(_19785_));
 sky130_fd_sc_hd__mux2_1 _23222_ (.A0(\cpuregs[1][18] ),
    .A1(_19785_),
    .S(_19784_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_2 _23223_ (.A(\cpuregs_wrdata[17] ),
    .X(_19786_));
 sky130_fd_sc_hd__mux2_1 _23224_ (.A0(\cpuregs[1][17] ),
    .A1(_19786_),
    .S(_19784_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_2 _23225_ (.A(\cpuregs_wrdata[16] ),
    .X(_19787_));
 sky130_fd_sc_hd__mux2_1 _23226_ (.A0(\cpuregs[1][16] ),
    .A1(_19787_),
    .S(_19784_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_2 _23227_ (.A(\cpuregs_wrdata[15] ),
    .X(_19788_));
 sky130_fd_sc_hd__mux2_1 _23228_ (.A0(\cpuregs[1][15] ),
    .A1(_19788_),
    .S(_19784_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_2 _23229_ (.A(\cpuregs_wrdata[14] ),
    .X(_19789_));
 sky130_fd_sc_hd__mux2_1 _23230_ (.A0(\cpuregs[1][14] ),
    .A1(_19789_),
    .S(_19784_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_2 _23231_ (.A(\cpuregs_wrdata[13] ),
    .X(_19790_));
 sky130_fd_sc_hd__buf_4 _23232_ (.A(_19769_),
    .X(_19791_));
 sky130_fd_sc_hd__mux2_1 _23233_ (.A0(\cpuregs[1][13] ),
    .A1(_19790_),
    .S(_19791_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_2 _23234_ (.A(\cpuregs_wrdata[12] ),
    .X(_19792_));
 sky130_fd_sc_hd__mux2_1 _23235_ (.A0(\cpuregs[1][12] ),
    .A1(_19792_),
    .S(_19791_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_2 _23236_ (.A(\cpuregs_wrdata[11] ),
    .X(_19793_));
 sky130_fd_sc_hd__mux2_1 _23237_ (.A0(\cpuregs[1][11] ),
    .A1(_19793_),
    .S(_19791_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_2 _23238_ (.A(\cpuregs_wrdata[10] ),
    .X(_19794_));
 sky130_fd_sc_hd__mux2_1 _23239_ (.A0(\cpuregs[1][10] ),
    .A1(_19794_),
    .S(_19791_),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_2 _23240_ (.A(\cpuregs_wrdata[9] ),
    .X(_19795_));
 sky130_fd_sc_hd__mux2_1 _23241_ (.A0(\cpuregs[1][9] ),
    .A1(_19795_),
    .S(_19791_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_2 _23242_ (.A(\cpuregs_wrdata[8] ),
    .X(_19796_));
 sky130_fd_sc_hd__mux2_1 _23243_ (.A0(\cpuregs[1][8] ),
    .A1(_19796_),
    .S(_19791_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_2 _23244_ (.A(\cpuregs_wrdata[7] ),
    .X(_19797_));
 sky130_fd_sc_hd__clkbuf_4 _23245_ (.A(_19768_),
    .X(_19798_));
 sky130_fd_sc_hd__mux2_1 _23246_ (.A0(\cpuregs[1][7] ),
    .A1(_19797_),
    .S(_19798_),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_2 _23247_ (.A(\cpuregs_wrdata[6] ),
    .X(_19799_));
 sky130_fd_sc_hd__mux2_1 _23248_ (.A0(\cpuregs[1][6] ),
    .A1(_19799_),
    .S(_19798_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_2 _23249_ (.A(\cpuregs_wrdata[5] ),
    .X(_19800_));
 sky130_fd_sc_hd__mux2_1 _23250_ (.A0(\cpuregs[1][5] ),
    .A1(_19800_),
    .S(_19798_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_2 _23251_ (.A(\cpuregs_wrdata[4] ),
    .X(_19801_));
 sky130_fd_sc_hd__mux2_1 _23252_ (.A0(\cpuregs[1][4] ),
    .A1(_19801_),
    .S(_19798_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_2 _23253_ (.A(\cpuregs_wrdata[3] ),
    .X(_19802_));
 sky130_fd_sc_hd__mux2_1 _23254_ (.A0(\cpuregs[1][3] ),
    .A1(_19802_),
    .S(_19798_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_2 _23255_ (.A(\cpuregs_wrdata[2] ),
    .X(_19803_));
 sky130_fd_sc_hd__mux2_1 _23256_ (.A0(\cpuregs[1][2] ),
    .A1(_19803_),
    .S(_19798_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_2 _23257_ (.A(\cpuregs_wrdata[1] ),
    .X(_19804_));
 sky130_fd_sc_hd__mux2_1 _23258_ (.A0(\cpuregs[1][1] ),
    .A1(_19804_),
    .S(_19769_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_2 _23259_ (.A(\cpuregs_wrdata[0] ),
    .X(_19805_));
 sky130_fd_sc_hd__mux2_1 _23260_ (.A0(\cpuregs[1][0] ),
    .A1(_19805_),
    .S(_19769_),
    .X(_03375_));
 sky130_fd_sc_hd__or3b_1 _23261_ (.A(_19592_),
    .B(_19599_),
    .C_N(_19712_),
    .X(_19806_));
 sky130_fd_sc_hd__buf_6 _23262_ (.A(_19806_),
    .X(_19807_));
 sky130_fd_sc_hd__clkbuf_4 _23263_ (.A(_19807_),
    .X(_19808_));
 sky130_fd_sc_hd__mux2_1 _23264_ (.A0(_19720_),
    .A1(\cpuregs[12][31] ),
    .S(_19808_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _23265_ (.A0(_19724_),
    .A1(\cpuregs[12][30] ),
    .S(_19808_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _23266_ (.A0(_19725_),
    .A1(\cpuregs[12][29] ),
    .S(_19808_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _23267_ (.A0(_19726_),
    .A1(\cpuregs[12][28] ),
    .S(_19808_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _23268_ (.A0(_19727_),
    .A1(\cpuregs[12][27] ),
    .S(_19808_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _23269_ (.A0(_19728_),
    .A1(\cpuregs[12][26] ),
    .S(_19808_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_4 _23270_ (.A(_19807_),
    .X(_19809_));
 sky130_fd_sc_hd__mux2_1 _23271_ (.A0(_19729_),
    .A1(\cpuregs[12][25] ),
    .S(_19809_),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_1 _23272_ (.A0(_19731_),
    .A1(\cpuregs[12][24] ),
    .S(_19809_),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _23273_ (.A0(_19732_),
    .A1(\cpuregs[12][23] ),
    .S(_19809_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _23274_ (.A0(_19733_),
    .A1(\cpuregs[12][22] ),
    .S(_19809_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_1 _23275_ (.A0(_19734_),
    .A1(\cpuregs[12][21] ),
    .S(_19809_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_1 _23276_ (.A0(_19735_),
    .A1(\cpuregs[12][20] ),
    .S(_19809_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_4 _23277_ (.A(_19807_),
    .X(_19810_));
 sky130_fd_sc_hd__mux2_1 _23278_ (.A0(_19736_),
    .A1(\cpuregs[12][19] ),
    .S(_19810_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_1 _23279_ (.A0(_19738_),
    .A1(\cpuregs[12][18] ),
    .S(_19810_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _23280_ (.A0(_19739_),
    .A1(\cpuregs[12][17] ),
    .S(_19810_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _23281_ (.A0(_19740_),
    .A1(\cpuregs[12][16] ),
    .S(_19810_),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_1 _23282_ (.A0(_19741_),
    .A1(\cpuregs[12][15] ),
    .S(_19810_),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _23283_ (.A0(_19742_),
    .A1(\cpuregs[12][14] ),
    .S(_19810_),
    .X(_03357_));
 sky130_fd_sc_hd__buf_4 _23284_ (.A(_19807_),
    .X(_19811_));
 sky130_fd_sc_hd__mux2_1 _23285_ (.A0(_19743_),
    .A1(\cpuregs[12][13] ),
    .S(_19811_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _23286_ (.A0(_19745_),
    .A1(\cpuregs[12][12] ),
    .S(_19811_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _23287_ (.A0(_19746_),
    .A1(\cpuregs[12][11] ),
    .S(_19811_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _23288_ (.A0(_19747_),
    .A1(\cpuregs[12][10] ),
    .S(_19811_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _23289_ (.A0(_19748_),
    .A1(\cpuregs[12][9] ),
    .S(_19811_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _23290_ (.A0(_19749_),
    .A1(\cpuregs[12][8] ),
    .S(_19811_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_4 _23291_ (.A(_19806_),
    .X(_19812_));
 sky130_fd_sc_hd__mux2_1 _23292_ (.A0(_19750_),
    .A1(\cpuregs[12][7] ),
    .S(_19812_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _23293_ (.A0(_19752_),
    .A1(\cpuregs[12][6] ),
    .S(_19812_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _23294_ (.A0(_19753_),
    .A1(\cpuregs[12][5] ),
    .S(_19812_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _23295_ (.A0(_19754_),
    .A1(\cpuregs[12][4] ),
    .S(_19812_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _23296_ (.A0(_19755_),
    .A1(\cpuregs[12][3] ),
    .S(_19812_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _23297_ (.A0(_19756_),
    .A1(\cpuregs[12][2] ),
    .S(_19812_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _23298_ (.A0(_19757_),
    .A1(\cpuregs[12][1] ),
    .S(_19807_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _23299_ (.A0(_19758_),
    .A1(\cpuregs[12][0] ),
    .S(_19807_),
    .X(_03343_));
 sky130_fd_sc_hd__or3_1 _23300_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C(_19592_),
    .X(_19813_));
 sky130_fd_sc_hd__nor2_1 _23301_ (.A(_19813_),
    .B(_19599_),
    .Y(_19814_));
 sky130_fd_sc_hd__buf_4 _23302_ (.A(_19814_),
    .X(_19815_));
 sky130_fd_sc_hd__clkbuf_4 _23303_ (.A(_19815_),
    .X(_19816_));
 sky130_fd_sc_hd__mux2_1 _23304_ (.A0(\cpuregs[16][31] ),
    .A1(_19767_),
    .S(_19816_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _23305_ (.A0(\cpuregs[16][30] ),
    .A1(_19771_),
    .S(_19816_),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_1 _23306_ (.A0(\cpuregs[16][29] ),
    .A1(_19772_),
    .S(_19816_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _23307_ (.A0(\cpuregs[16][28] ),
    .A1(_19773_),
    .S(_19816_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _23308_ (.A0(\cpuregs[16][27] ),
    .A1(_19774_),
    .S(_19816_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _23309_ (.A0(\cpuregs[16][26] ),
    .A1(_19775_),
    .S(_19816_),
    .X(_03337_));
 sky130_fd_sc_hd__buf_4 _23310_ (.A(_19815_),
    .X(_19817_));
 sky130_fd_sc_hd__mux2_1 _23311_ (.A0(\cpuregs[16][25] ),
    .A1(_19776_),
    .S(_19817_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_1 _23312_ (.A0(\cpuregs[16][24] ),
    .A1(_19778_),
    .S(_19817_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _23313_ (.A0(\cpuregs[16][23] ),
    .A1(_19779_),
    .S(_19817_),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _23314_ (.A0(\cpuregs[16][22] ),
    .A1(_19780_),
    .S(_19817_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _23315_ (.A0(\cpuregs[16][21] ),
    .A1(_19781_),
    .S(_19817_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _23316_ (.A0(\cpuregs[16][20] ),
    .A1(_19782_),
    .S(_19817_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_4 _23317_ (.A(_19815_),
    .X(_19818_));
 sky130_fd_sc_hd__mux2_1 _23318_ (.A0(\cpuregs[16][19] ),
    .A1(_19783_),
    .S(_19818_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _23319_ (.A0(\cpuregs[16][18] ),
    .A1(_19785_),
    .S(_19818_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _23320_ (.A0(\cpuregs[16][17] ),
    .A1(_19786_),
    .S(_19818_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _23321_ (.A0(\cpuregs[16][16] ),
    .A1(_19787_),
    .S(_19818_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _23322_ (.A0(\cpuregs[16][15] ),
    .A1(_19788_),
    .S(_19818_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_1 _23323_ (.A0(\cpuregs[16][14] ),
    .A1(_19789_),
    .S(_19818_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_4 _23324_ (.A(_19815_),
    .X(_19819_));
 sky130_fd_sc_hd__mux2_1 _23325_ (.A0(\cpuregs[16][13] ),
    .A1(_19790_),
    .S(_19819_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _23326_ (.A0(\cpuregs[16][12] ),
    .A1(_19792_),
    .S(_19819_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _23327_ (.A0(\cpuregs[16][11] ),
    .A1(_19793_),
    .S(_19819_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_1 _23328_ (.A0(\cpuregs[16][10] ),
    .A1(_19794_),
    .S(_19819_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_1 _23329_ (.A0(\cpuregs[16][9] ),
    .A1(_19795_),
    .S(_19819_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _23330_ (.A0(\cpuregs[16][8] ),
    .A1(_19796_),
    .S(_19819_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_4 _23331_ (.A(_19814_),
    .X(_19820_));
 sky130_fd_sc_hd__mux2_1 _23332_ (.A0(\cpuregs[16][7] ),
    .A1(_19797_),
    .S(_19820_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _23333_ (.A0(\cpuregs[16][6] ),
    .A1(_19799_),
    .S(_19820_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_1 _23334_ (.A0(\cpuregs[16][5] ),
    .A1(_19800_),
    .S(_19820_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_1 _23335_ (.A0(\cpuregs[16][4] ),
    .A1(_19801_),
    .S(_19820_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _23336_ (.A0(\cpuregs[16][3] ),
    .A1(_19802_),
    .S(_19820_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _23337_ (.A0(\cpuregs[16][2] ),
    .A1(_19803_),
    .S(_19820_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_1 _23338_ (.A0(\cpuregs[16][1] ),
    .A1(_19804_),
    .S(_19815_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_1 _23339_ (.A0(\cpuregs[16][0] ),
    .A1(_19805_),
    .S(_19815_),
    .X(_03311_));
 sky130_fd_sc_hd__and2_1 _23340_ (.A(_19642_),
    .B(_19687_),
    .X(_19821_));
 sky130_fd_sc_hd__buf_4 _23341_ (.A(_19821_),
    .X(_19822_));
 sky130_fd_sc_hd__clkbuf_4 _23342_ (.A(_19822_),
    .X(_19823_));
 sky130_fd_sc_hd__mux2_1 _23343_ (.A0(\cpuregs[17][31] ),
    .A1(_19767_),
    .S(_19823_),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_1 _23344_ (.A0(\cpuregs[17][30] ),
    .A1(_19771_),
    .S(_19823_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _23345_ (.A0(\cpuregs[17][29] ),
    .A1(_19772_),
    .S(_19823_),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_1 _23346_ (.A0(\cpuregs[17][28] ),
    .A1(_19773_),
    .S(_19823_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _23347_ (.A0(\cpuregs[17][27] ),
    .A1(_19774_),
    .S(_19823_),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _23348_ (.A0(\cpuregs[17][26] ),
    .A1(_19775_),
    .S(_19823_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_4 _23349_ (.A(_19822_),
    .X(_19824_));
 sky130_fd_sc_hd__mux2_1 _23350_ (.A0(\cpuregs[17][25] ),
    .A1(_19776_),
    .S(_19824_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_1 _23351_ (.A0(\cpuregs[17][24] ),
    .A1(_19778_),
    .S(_19824_),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_1 _23352_ (.A0(\cpuregs[17][23] ),
    .A1(_19779_),
    .S(_19824_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _23353_ (.A0(\cpuregs[17][22] ),
    .A1(_19780_),
    .S(_19824_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _23354_ (.A0(\cpuregs[17][21] ),
    .A1(_19781_),
    .S(_19824_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _23355_ (.A0(\cpuregs[17][20] ),
    .A1(_19782_),
    .S(_19824_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_4 _23356_ (.A(_19822_),
    .X(_19825_));
 sky130_fd_sc_hd__mux2_1 _23357_ (.A0(\cpuregs[17][19] ),
    .A1(_19783_),
    .S(_19825_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _23358_ (.A0(\cpuregs[17][18] ),
    .A1(_19785_),
    .S(_19825_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _23359_ (.A0(\cpuregs[17][17] ),
    .A1(_19786_),
    .S(_19825_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _23360_ (.A0(\cpuregs[17][16] ),
    .A1(_19787_),
    .S(_19825_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _23361_ (.A0(\cpuregs[17][15] ),
    .A1(_19788_),
    .S(_19825_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _23362_ (.A0(\cpuregs[17][14] ),
    .A1(_19789_),
    .S(_19825_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_4 _23363_ (.A(_19822_),
    .X(_19826_));
 sky130_fd_sc_hd__mux2_1 _23364_ (.A0(\cpuregs[17][13] ),
    .A1(_19790_),
    .S(_19826_),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _23365_ (.A0(\cpuregs[17][12] ),
    .A1(_19792_),
    .S(_19826_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _23366_ (.A0(\cpuregs[17][11] ),
    .A1(_19793_),
    .S(_19826_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _23367_ (.A0(\cpuregs[17][10] ),
    .A1(_19794_),
    .S(_19826_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _23368_ (.A0(\cpuregs[17][9] ),
    .A1(_19795_),
    .S(_19826_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _23369_ (.A0(\cpuregs[17][8] ),
    .A1(_19796_),
    .S(_19826_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_4 _23370_ (.A(_19821_),
    .X(_19827_));
 sky130_fd_sc_hd__mux2_1 _23371_ (.A0(\cpuregs[17][7] ),
    .A1(_19797_),
    .S(_19827_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _23372_ (.A0(\cpuregs[17][6] ),
    .A1(_19799_),
    .S(_19827_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _23373_ (.A0(\cpuregs[17][5] ),
    .A1(_19800_),
    .S(_19827_),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _23374_ (.A0(\cpuregs[17][4] ),
    .A1(_19801_),
    .S(_19827_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _23375_ (.A0(\cpuregs[17][3] ),
    .A1(_19802_),
    .S(_19827_),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_1 _23376_ (.A0(\cpuregs[17][2] ),
    .A1(_19803_),
    .S(_19827_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_1 _23377_ (.A0(\cpuregs[17][1] ),
    .A1(_19804_),
    .S(_19822_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _23378_ (.A0(\cpuregs[17][0] ),
    .A1(_19805_),
    .S(_19822_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_4 _23379_ (.A(\pcpi_mul.rs2[31] ),
    .X(_19828_));
 sky130_fd_sc_hd__buf_8 _23380_ (.A(_19828_),
    .X(_19829_));
 sky130_fd_sc_hd__clkbuf_2 _23381_ (.A(_19829_),
    .X(_19830_));
 sky130_fd_sc_hd__clkbuf_2 _23382_ (.A(_19830_),
    .X(_19831_));
 sky130_fd_sc_hd__a21o_1 _23383_ (.A1(_19831_),
    .A2(_18689_),
    .B1(_18691_),
    .X(_03278_));
 sky130_fd_sc_hd__buf_4 _23384_ (.A(\pcpi_mul.rs2[30] ),
    .X(_19832_));
 sky130_fd_sc_hd__buf_4 _23385_ (.A(_19832_),
    .X(_19833_));
 sky130_fd_sc_hd__buf_2 _23386_ (.A(_19833_),
    .X(_19834_));
 sky130_fd_sc_hd__mux2_1 _23387_ (.A0(net361),
    .A1(_19834_),
    .S(_18689_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_6 _23388_ (.A(\pcpi_mul.rs2[29] ),
    .X(_19835_));
 sky130_fd_sc_hd__buf_4 _23389_ (.A(_19835_),
    .X(_19836_));
 sky130_fd_sc_hd__buf_2 _23390_ (.A(_19836_),
    .X(_19837_));
 sky130_fd_sc_hd__buf_2 _23391_ (.A(_18680_),
    .X(_19838_));
 sky130_fd_sc_hd__mux2_1 _23392_ (.A0(_19655_),
    .A1(_19837_),
    .S(_19838_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_4 _23393_ (.A(\pcpi_mul.rs2[28] ),
    .X(_19839_));
 sky130_fd_sc_hd__buf_6 _23394_ (.A(_19839_),
    .X(_19840_));
 sky130_fd_sc_hd__buf_6 _23395_ (.A(_19840_),
    .X(_19841_));
 sky130_fd_sc_hd__buf_2 _23396_ (.A(_19841_),
    .X(_19842_));
 sky130_fd_sc_hd__mux2_1 _23397_ (.A0(net358),
    .A1(_19842_),
    .S(_19838_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_6 _23398_ (.A(\pcpi_mul.rs2[27] ),
    .X(_19843_));
 sky130_fd_sc_hd__buf_4 _23399_ (.A(_19843_),
    .X(_19844_));
 sky130_fd_sc_hd__clkbuf_4 _23400_ (.A(_19844_),
    .X(_19845_));
 sky130_fd_sc_hd__mux2_1 _23401_ (.A0(_19656_),
    .A1(_19845_),
    .S(_19838_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_4 _23402_ (.A(\pcpi_mul.rs2[26] ),
    .X(_19846_));
 sky130_fd_sc_hd__buf_6 _23403_ (.A(_19846_),
    .X(_19847_));
 sky130_fd_sc_hd__buf_6 _23404_ (.A(_19847_),
    .X(_19848_));
 sky130_fd_sc_hd__clkbuf_4 _23405_ (.A(_19848_),
    .X(_19849_));
 sky130_fd_sc_hd__mux2_1 _23406_ (.A0(_19657_),
    .A1(_19849_),
    .S(_19838_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_4 _23407_ (.A(\pcpi_mul.rs2[25] ),
    .X(_19850_));
 sky130_fd_sc_hd__buf_6 _23408_ (.A(_19850_),
    .X(_19851_));
 sky130_fd_sc_hd__buf_6 _23409_ (.A(_19851_),
    .X(_19852_));
 sky130_fd_sc_hd__mux2_1 _23410_ (.A0(_19659_),
    .A1(_19852_),
    .S(_19838_),
    .X(_03272_));
 sky130_fd_sc_hd__buf_2 _23411_ (.A(\pcpi_mul.rs2[24] ),
    .X(_19853_));
 sky130_fd_sc_hd__buf_6 _23412_ (.A(_19853_),
    .X(_19854_));
 sky130_fd_sc_hd__clkbuf_4 _23413_ (.A(_19854_),
    .X(_19855_));
 sky130_fd_sc_hd__clkbuf_4 _23414_ (.A(_19855_),
    .X(_19856_));
 sky130_fd_sc_hd__mux2_1 _23415_ (.A0(net354),
    .A1(_19856_),
    .S(_19838_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_4 _23416_ (.A(\pcpi_mul.rs2[23] ),
    .X(_19857_));
 sky130_fd_sc_hd__clkbuf_4 _23417_ (.A(_19857_),
    .X(_19858_));
 sky130_fd_sc_hd__buf_4 _23418_ (.A(_19858_),
    .X(_19859_));
 sky130_fd_sc_hd__buf_4 _23419_ (.A(_19859_),
    .X(_19860_));
 sky130_fd_sc_hd__buf_2 _23420_ (.A(_18680_),
    .X(_19861_));
 sky130_fd_sc_hd__mux2_1 _23421_ (.A0(net353),
    .A1(_19860_),
    .S(_19861_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_4 _23422_ (.A(\pcpi_mul.rs2[22] ),
    .X(_19862_));
 sky130_fd_sc_hd__buf_6 _23423_ (.A(_19862_),
    .X(_19863_));
 sky130_fd_sc_hd__buf_4 _23424_ (.A(_19863_),
    .X(_19864_));
 sky130_fd_sc_hd__mux2_1 _23425_ (.A0(net352),
    .A1(_19864_),
    .S(_19861_),
    .X(_03269_));
 sky130_fd_sc_hd__buf_6 _23426_ (.A(\pcpi_mul.rs2[21] ),
    .X(_19865_));
 sky130_fd_sc_hd__clkbuf_8 _23427_ (.A(_19865_),
    .X(_19866_));
 sky130_fd_sc_hd__clkbuf_4 _23428_ (.A(_19866_),
    .X(_19867_));
 sky130_fd_sc_hd__buf_4 _23429_ (.A(_19867_),
    .X(_19868_));
 sky130_fd_sc_hd__mux2_1 _23430_ (.A0(_19660_),
    .A1(_19868_),
    .S(_19861_),
    .X(_03268_));
 sky130_fd_sc_hd__clkbuf_4 _23431_ (.A(\pcpi_mul.rs2[20] ),
    .X(_19869_));
 sky130_fd_sc_hd__buf_6 _23432_ (.A(_19869_),
    .X(_19870_));
 sky130_fd_sc_hd__buf_4 _23433_ (.A(_19870_),
    .X(_19871_));
 sky130_fd_sc_hd__mux2_1 _23434_ (.A0(net350),
    .A1(_19871_),
    .S(_19861_),
    .X(_03267_));
 sky130_fd_sc_hd__clkbuf_4 _23435_ (.A(\pcpi_mul.rs2[19] ),
    .X(_19872_));
 sky130_fd_sc_hd__buf_6 _23436_ (.A(_19872_),
    .X(_19873_));
 sky130_fd_sc_hd__buf_8 _23437_ (.A(_19873_),
    .X(_19874_));
 sky130_fd_sc_hd__buf_6 _23438_ (.A(_19874_),
    .X(_19875_));
 sky130_fd_sc_hd__mux2_1 _23439_ (.A0(net348),
    .A1(_19875_),
    .S(_19861_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_4 _23440_ (.A(\pcpi_mul.rs2[18] ),
    .X(_19876_));
 sky130_fd_sc_hd__clkbuf_4 _23441_ (.A(_19876_),
    .X(_19877_));
 sky130_fd_sc_hd__clkbuf_2 _23442_ (.A(_19877_),
    .X(_19878_));
 sky130_fd_sc_hd__buf_6 _23443_ (.A(net457),
    .X(_19879_));
 sky130_fd_sc_hd__mux2_1 _23444_ (.A0(_19662_),
    .A1(_19879_),
    .S(_19861_),
    .X(_03265_));
 sky130_fd_sc_hd__buf_4 _23445_ (.A(\pcpi_mul.rs2[17] ),
    .X(_19880_));
 sky130_fd_sc_hd__buf_6 _23446_ (.A(_19880_),
    .X(_19881_));
 sky130_fd_sc_hd__buf_6 _23447_ (.A(_19881_),
    .X(_19882_));
 sky130_fd_sc_hd__clkbuf_4 _23448_ (.A(_18679_),
    .X(_19883_));
 sky130_fd_sc_hd__clkbuf_4 _23449_ (.A(_19883_),
    .X(_19884_));
 sky130_fd_sc_hd__mux2_1 _23450_ (.A0(_19663_),
    .A1(_19882_),
    .S(_19884_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_2 _23451_ (.A(\pcpi_mul.rs2[16] ),
    .X(_19885_));
 sky130_fd_sc_hd__buf_4 _23452_ (.A(_19885_),
    .X(_19886_));
 sky130_fd_sc_hd__buf_4 _23453_ (.A(_19886_),
    .X(_19887_));
 sky130_fd_sc_hd__buf_4 _23454_ (.A(_19887_),
    .X(_19888_));
 sky130_fd_sc_hd__mux2_1 _23455_ (.A0(net345),
    .A1(_19888_),
    .S(_19884_),
    .X(_03263_));
 sky130_fd_sc_hd__buf_6 _23456_ (.A(\pcpi_mul.rs2[15] ),
    .X(_19889_));
 sky130_fd_sc_hd__buf_6 _23457_ (.A(_19889_),
    .X(_19890_));
 sky130_fd_sc_hd__clkbuf_2 _23458_ (.A(_19890_),
    .X(_19891_));
 sky130_fd_sc_hd__mux2_1 _23459_ (.A0(_19664_),
    .A1(_19891_),
    .S(_19884_),
    .X(_03262_));
 sky130_fd_sc_hd__buf_6 _23460_ (.A(\pcpi_mul.rs2[14] ),
    .X(_19892_));
 sky130_fd_sc_hd__buf_6 _23461_ (.A(_19892_),
    .X(_19893_));
 sky130_fd_sc_hd__buf_6 _23462_ (.A(_19893_),
    .X(_19894_));
 sky130_fd_sc_hd__mux2_1 _23463_ (.A0(net343),
    .A1(_19894_),
    .S(_19884_),
    .X(_03261_));
 sky130_fd_sc_hd__clkbuf_4 _23464_ (.A(\pcpi_mul.rs2[13] ),
    .X(_19895_));
 sky130_fd_sc_hd__buf_6 _23465_ (.A(_19895_),
    .X(_19896_));
 sky130_fd_sc_hd__buf_6 _23466_ (.A(_19896_),
    .X(_19897_));
 sky130_fd_sc_hd__mux2_1 _23467_ (.A0(_19666_),
    .A1(_19897_),
    .S(_19884_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_6 _23468_ (.A(\pcpi_mul.rs2[12] ),
    .X(_19898_));
 sky130_fd_sc_hd__buf_6 _23469_ (.A(_19898_),
    .X(_19899_));
 sky130_fd_sc_hd__buf_1 _23470_ (.A(_19899_),
    .X(_19900_));
 sky130_fd_sc_hd__mux2_1 _23471_ (.A0(net341),
    .A1(net455),
    .S(_19884_),
    .X(_03259_));
 sky130_fd_sc_hd__buf_6 _23472_ (.A(\pcpi_mul.rs2[11] ),
    .X(_19901_));
 sky130_fd_sc_hd__buf_6 _23473_ (.A(_19901_),
    .X(_19902_));
 sky130_fd_sc_hd__buf_6 _23474_ (.A(_19902_),
    .X(_19903_));
 sky130_fd_sc_hd__clkbuf_4 _23475_ (.A(_19883_),
    .X(_19904_));
 sky130_fd_sc_hd__mux2_1 _23476_ (.A0(_19667_),
    .A1(_19903_),
    .S(_19904_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_6 _23477_ (.A(\pcpi_mul.rs2[10] ),
    .X(_19905_));
 sky130_fd_sc_hd__buf_6 _23478_ (.A(_19905_),
    .X(_19906_));
 sky130_fd_sc_hd__buf_6 _23479_ (.A(_19906_),
    .X(_19907_));
 sky130_fd_sc_hd__mux2_1 _23480_ (.A0(net339),
    .A1(_19907_),
    .S(_19904_),
    .X(_03257_));
 sky130_fd_sc_hd__buf_6 _23481_ (.A(\pcpi_mul.rs2[9] ),
    .X(_19908_));
 sky130_fd_sc_hd__buf_6 _23482_ (.A(_19908_),
    .X(_19909_));
 sky130_fd_sc_hd__clkbuf_8 _23483_ (.A(_19909_),
    .X(_19910_));
 sky130_fd_sc_hd__mux2_1 _23484_ (.A0(_19668_),
    .A1(_19910_),
    .S(_19904_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_6 _23485_ (.A(\pcpi_mul.rs2[8] ),
    .X(_19911_));
 sky130_fd_sc_hd__buf_8 _23486_ (.A(_19911_),
    .X(_19912_));
 sky130_fd_sc_hd__buf_4 _23487_ (.A(_19912_),
    .X(_19913_));
 sky130_fd_sc_hd__mux2_1 _23488_ (.A0(net368),
    .A1(_19913_),
    .S(_19904_),
    .X(_03255_));
 sky130_fd_sc_hd__buf_6 _23489_ (.A(\pcpi_mul.rs2[7] ),
    .X(_19914_));
 sky130_fd_sc_hd__clkbuf_8 _23490_ (.A(_19914_),
    .X(_19915_));
 sky130_fd_sc_hd__buf_6 _23491_ (.A(_19915_),
    .X(_19916_));
 sky130_fd_sc_hd__mux2_1 _23492_ (.A0(_19670_),
    .A1(_19916_),
    .S(_19904_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_4 _23493_ (.A(\pcpi_mul.rs2[6] ),
    .X(_19917_));
 sky130_fd_sc_hd__buf_8 _23494_ (.A(_19917_),
    .X(_19918_));
 sky130_fd_sc_hd__mux2_1 _23495_ (.A0(_19671_),
    .A1(_19918_),
    .S(_19904_),
    .X(_03253_));
 sky130_fd_sc_hd__clkbuf_8 _23496_ (.A(\pcpi_mul.rs2[5] ),
    .X(_19919_));
 sky130_fd_sc_hd__buf_6 _23497_ (.A(_19919_),
    .X(_19920_));
 sky130_fd_sc_hd__clkbuf_4 _23498_ (.A(_19920_),
    .X(_19921_));
 sky130_fd_sc_hd__clkbuf_4 _23499_ (.A(_19883_),
    .X(_19922_));
 sky130_fd_sc_hd__mux2_1 _23500_ (.A0(_19672_),
    .A1(_19921_),
    .S(_19922_),
    .X(_03252_));
 sky130_fd_sc_hd__clkbuf_4 _23501_ (.A(\pcpi_mul.rs2[4] ),
    .X(_19923_));
 sky130_fd_sc_hd__buf_4 _23502_ (.A(_19923_),
    .X(_19924_));
 sky130_fd_sc_hd__buf_6 _23503_ (.A(_19924_),
    .X(_19925_));
 sky130_fd_sc_hd__buf_4 _23504_ (.A(_19925_),
    .X(_19926_));
 sky130_fd_sc_hd__mux2_1 _23505_ (.A0(_19673_),
    .A1(_19926_),
    .S(_19922_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_4 _23506_ (.A(\pcpi_mul.rs2[3] ),
    .X(_19927_));
 sky130_fd_sc_hd__buf_8 _23507_ (.A(_19927_),
    .X(_19928_));
 sky130_fd_sc_hd__buf_6 _23508_ (.A(_19928_),
    .X(_19929_));
 sky130_fd_sc_hd__mux2_1 _23509_ (.A0(_19674_),
    .A1(_19929_),
    .S(_19922_),
    .X(_03250_));
 sky130_fd_sc_hd__buf_2 _23510_ (.A(\pcpi_mul.rs2[2] ),
    .X(_19930_));
 sky130_fd_sc_hd__buf_6 _23511_ (.A(_19930_),
    .X(_19931_));
 sky130_fd_sc_hd__buf_4 _23512_ (.A(_19931_),
    .X(_19932_));
 sky130_fd_sc_hd__mux2_1 _23513_ (.A0(_19675_),
    .A1(_19932_),
    .S(_19922_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_4 _23514_ (.A(\pcpi_mul.rs2[1] ),
    .X(_19933_));
 sky130_fd_sc_hd__clkbuf_4 _23515_ (.A(_19933_),
    .X(_19934_));
 sky130_fd_sc_hd__buf_4 _23516_ (.A(_19934_),
    .X(_19935_));
 sky130_fd_sc_hd__mux2_1 _23517_ (.A0(_19676_),
    .A1(_19935_),
    .S(_19922_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_4 _23518_ (.A(\pcpi_mul.rs2[0] ),
    .X(_19936_));
 sky130_fd_sc_hd__buf_8 _23519_ (.A(_19936_),
    .X(_19937_));
 sky130_fd_sc_hd__buf_6 _23520_ (.A(_19937_),
    .X(_19938_));
 sky130_fd_sc_hd__clkbuf_8 _23521_ (.A(_19938_),
    .X(_19939_));
 sky130_fd_sc_hd__mux2_1 _23522_ (.A0(_19677_),
    .A1(_19939_),
    .S(_19922_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _23523_ (.A0(net273),
    .A1(_02541_),
    .S(_18569_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _23524_ (.A0(net272),
    .A1(_02540_),
    .S(_18569_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _23525_ (.A0(net271),
    .A1(_02539_),
    .S(_18568_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_1 _23526_ (.A0(net270),
    .A1(_02538_),
    .S(_18568_),
    .X(_03243_));
 sky130_vsdinv _23527_ (.A(_00330_),
    .Y(_19940_));
 sky130_fd_sc_hd__and4_1 _23528_ (.A(_18577_),
    .B(_18579_),
    .C(_19940_),
    .D(_18581_),
    .X(_19941_));
 sky130_fd_sc_hd__clkbuf_2 _23529_ (.A(_18860_),
    .X(_19942_));
 sky130_fd_sc_hd__a32o_1 _23530_ (.A1(_19941_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(is_alu_reg_reg),
    .B2(_19942_),
    .X(_03242_));
 sky130_vsdinv _23531_ (.A(_00329_),
    .Y(_19943_));
 sky130_fd_sc_hd__a32o_1 _23532_ (.A1(_19941_),
    .A2(_19943_),
    .A3(_00328_),
    .B1(is_alu_reg_imm),
    .B2(_19942_),
    .X(_03241_));
 sky130_fd_sc_hd__and2_1 _23533_ (.A(_19642_),
    .B(_19712_),
    .X(_19944_));
 sky130_fd_sc_hd__buf_6 _23534_ (.A(_19944_),
    .X(_19945_));
 sky130_fd_sc_hd__clkbuf_4 _23535_ (.A(_19945_),
    .X(_19946_));
 sky130_fd_sc_hd__mux2_1 _23536_ (.A0(\cpuregs[13][31] ),
    .A1(\cpuregs_wrdata[31] ),
    .S(_19946_),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _23537_ (.A0(\cpuregs[13][30] ),
    .A1(\cpuregs_wrdata[30] ),
    .S(_19946_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _23538_ (.A0(\cpuregs[13][29] ),
    .A1(\cpuregs_wrdata[29] ),
    .S(_19946_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _23539_ (.A0(\cpuregs[13][28] ),
    .A1(\cpuregs_wrdata[28] ),
    .S(_19946_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _23540_ (.A0(\cpuregs[13][27] ),
    .A1(\cpuregs_wrdata[27] ),
    .S(_19946_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_1 _23541_ (.A0(\cpuregs[13][26] ),
    .A1(\cpuregs_wrdata[26] ),
    .S(_19946_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_4 _23542_ (.A(_19945_),
    .X(_19947_));
 sky130_fd_sc_hd__mux2_1 _23543_ (.A0(\cpuregs[13][25] ),
    .A1(\cpuregs_wrdata[25] ),
    .S(_19947_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _23544_ (.A0(\cpuregs[13][24] ),
    .A1(\cpuregs_wrdata[24] ),
    .S(_19947_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _23545_ (.A0(\cpuregs[13][23] ),
    .A1(\cpuregs_wrdata[23] ),
    .S(_19947_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _23546_ (.A0(\cpuregs[13][22] ),
    .A1(\cpuregs_wrdata[22] ),
    .S(_19947_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _23547_ (.A0(\cpuregs[13][21] ),
    .A1(\cpuregs_wrdata[21] ),
    .S(_19947_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _23548_ (.A0(\cpuregs[13][20] ),
    .A1(\cpuregs_wrdata[20] ),
    .S(_19947_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_4 _23549_ (.A(_19945_),
    .X(_19948_));
 sky130_fd_sc_hd__mux2_1 _23550_ (.A0(\cpuregs[13][19] ),
    .A1(\cpuregs_wrdata[19] ),
    .S(_19948_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_1 _23551_ (.A0(\cpuregs[13][18] ),
    .A1(\cpuregs_wrdata[18] ),
    .S(_19948_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _23552_ (.A0(\cpuregs[13][17] ),
    .A1(\cpuregs_wrdata[17] ),
    .S(_19948_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _23553_ (.A0(\cpuregs[13][16] ),
    .A1(\cpuregs_wrdata[16] ),
    .S(_19948_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _23554_ (.A0(\cpuregs[13][15] ),
    .A1(\cpuregs_wrdata[15] ),
    .S(_19948_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _23555_ (.A0(\cpuregs[13][14] ),
    .A1(\cpuregs_wrdata[14] ),
    .S(_19948_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_4 _23556_ (.A(_19945_),
    .X(_19949_));
 sky130_fd_sc_hd__mux2_1 _23557_ (.A0(\cpuregs[13][13] ),
    .A1(\cpuregs_wrdata[13] ),
    .S(_19949_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _23558_ (.A0(\cpuregs[13][12] ),
    .A1(\cpuregs_wrdata[12] ),
    .S(_19949_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _23559_ (.A0(\cpuregs[13][11] ),
    .A1(\cpuregs_wrdata[11] ),
    .S(_19949_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_1 _23560_ (.A0(\cpuregs[13][10] ),
    .A1(\cpuregs_wrdata[10] ),
    .S(_19949_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _23561_ (.A0(\cpuregs[13][9] ),
    .A1(\cpuregs_wrdata[9] ),
    .S(_19949_),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _23562_ (.A0(\cpuregs[13][8] ),
    .A1(\cpuregs_wrdata[8] ),
    .S(_19949_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_2 _23563_ (.A(_19944_),
    .X(_19950_));
 sky130_fd_sc_hd__mux2_1 _23564_ (.A0(\cpuregs[13][7] ),
    .A1(\cpuregs_wrdata[7] ),
    .S(_19950_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _23565_ (.A0(\cpuregs[13][6] ),
    .A1(\cpuregs_wrdata[6] ),
    .S(_19950_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_1 _23566_ (.A0(\cpuregs[13][5] ),
    .A1(\cpuregs_wrdata[5] ),
    .S(_19950_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_1 _23567_ (.A0(\cpuregs[13][4] ),
    .A1(\cpuregs_wrdata[4] ),
    .S(_19950_),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_1 _23568_ (.A0(\cpuregs[13][3] ),
    .A1(\cpuregs_wrdata[3] ),
    .S(_19950_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_1 _23569_ (.A0(\cpuregs[13][2] ),
    .A1(\cpuregs_wrdata[2] ),
    .S(_19950_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _23570_ (.A0(\cpuregs[13][1] ),
    .A1(\cpuregs_wrdata[1] ),
    .S(_19945_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _23571_ (.A0(\cpuregs[13][0] ),
    .A1(\cpuregs_wrdata[0] ),
    .S(_19945_),
    .X(_03209_));
 sky130_fd_sc_hd__buf_2 _23572_ (.A(is_sb_sh_sw),
    .X(_19951_));
 sky130_fd_sc_hd__a32o_1 _23573_ (.A1(_19941_),
    .A2(_00329_),
    .A3(_18858_),
    .B1(_19951_),
    .B2(_19942_),
    .X(_03208_));
 sky130_fd_sc_hd__nor2_1 _23574_ (.A(instr_jalr),
    .B(_18905_),
    .Y(_19952_));
 sky130_fd_sc_hd__a31o_1 _23575_ (.A1(_18915_),
    .A2(_18919_),
    .A3(_00335_),
    .B1(_18932_),
    .X(_19953_));
 sky130_fd_sc_hd__clkbuf_2 _23576_ (.A(_18917_),
    .X(_19954_));
 sky130_fd_sc_hd__clkbuf_4 _23577_ (.A(_19954_),
    .X(_19955_));
 sky130_fd_sc_hd__o2bb2a_1 _23578_ (.A1_N(_19952_),
    .A2_N(_19953_),
    .B1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B2(_19955_),
    .X(_03207_));
 sky130_fd_sc_hd__and3_1 _23579_ (.A(_18885_),
    .B(_18876_),
    .C(_18880_),
    .X(_19956_));
 sky130_fd_sc_hd__o2111a_1 _23580_ (.A1(_18893_),
    .A2(_18877_),
    .B1(_18878_),
    .C1(_18873_),
    .D1(_18889_),
    .X(_19957_));
 sky130_fd_sc_hd__buf_6 _23581_ (.A(is_slli_srli_srai),
    .X(_19958_));
 sky130_fd_sc_hd__clkbuf_2 _23582_ (.A(_18930_),
    .X(_19959_));
 sky130_fd_sc_hd__a32o_1 _23583_ (.A1(_19956_),
    .A2(_18933_),
    .A3(_19957_),
    .B1(_19958_),
    .B2(_19959_),
    .X(_03206_));
 sky130_fd_sc_hd__a32o_1 _23584_ (.A1(_19941_),
    .A2(_19943_),
    .A3(_18858_),
    .B1(is_lb_lh_lw_lbu_lhu),
    .B2(_19942_),
    .X(_03205_));
 sky130_fd_sc_hd__buf_4 _23585_ (.A(\decoded_imm_uj[20] ),
    .X(_19960_));
 sky130_fd_sc_hd__buf_6 _23586_ (.A(_19960_),
    .X(_19961_));
 sky130_fd_sc_hd__buf_4 _23587_ (.A(_19961_),
    .X(_19962_));
 sky130_fd_sc_hd__mux2_4 _23588_ (.A0(_19962_),
    .A1(\mem_rdata_latched[31] ),
    .S(_18862_),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_1 _23589_ (.A0(\decoded_imm_uj[19] ),
    .A1(\mem_rdata_latched[19] ),
    .S(_18862_),
    .X(_03203_));
 sky130_vsdinv _23590_ (.A(\decoded_imm_uj[18] ),
    .Y(_19963_));
 sky130_fd_sc_hd__o21ai_1 _23591_ (.A1(_19963_),
    .A2(_21108_),
    .B1(_18863_),
    .Y(_03202_));
 sky130_vsdinv _23592_ (.A(\decoded_imm_uj[17] ),
    .Y(_19964_));
 sky130_fd_sc_hd__o21ai_1 _23593_ (.A1(_19964_),
    .A2(_21108_),
    .B1(_18864_),
    .Y(_03201_));
 sky130_vsdinv _23594_ (.A(\decoded_imm_uj[16] ),
    .Y(_19965_));
 sky130_fd_sc_hd__o21ai_1 _23595_ (.A1(_19965_),
    .A2(_21108_),
    .B1(_18865_),
    .Y(_03200_));
 sky130_vsdinv _23596_ (.A(\decoded_imm_uj[15] ),
    .Y(_19966_));
 sky130_fd_sc_hd__o21ai_1 _23597_ (.A1(_19966_),
    .A2(_21108_),
    .B1(_18866_),
    .Y(_03199_));
 sky130_fd_sc_hd__buf_2 _23598_ (.A(_18577_),
    .X(_19967_));
 sky130_fd_sc_hd__mux2_1 _23599_ (.A0(\decoded_imm_uj[14] ),
    .A1(\mem_rdata_latched[14] ),
    .S(_19967_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_1 _23600_ (.A0(\decoded_imm_uj[13] ),
    .A1(\mem_rdata_latched[13] ),
    .S(_19967_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_1 _23601_ (.A0(\decoded_imm_uj[12] ),
    .A1(\mem_rdata_latched[12] ),
    .S(_19967_),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_1 _23602_ (.A0(\decoded_imm_uj[11] ),
    .A1(\mem_rdata_latched[20] ),
    .S(_19967_),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_1 _23603_ (.A0(\decoded_imm_uj[10] ),
    .A1(\mem_rdata_latched[30] ),
    .S(_19967_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _23604_ (.A0(\decoded_imm_uj[9] ),
    .A1(\mem_rdata_latched[29] ),
    .S(_19967_),
    .X(_03193_));
 sky130_fd_sc_hd__buf_2 _23605_ (.A(_18577_),
    .X(_19968_));
 sky130_fd_sc_hd__mux2_1 _23606_ (.A0(\decoded_imm_uj[8] ),
    .A1(\mem_rdata_latched[28] ),
    .S(_19968_),
    .X(_03192_));
 sky130_fd_sc_hd__and3_1 _23607_ (.A(_18573_),
    .B(mem_do_rinst),
    .C(\mem_rdata_latched[27] ),
    .X(_19969_));
 sky130_fd_sc_hd__a21o_1 _23608_ (.A1(_00337_),
    .A2(\decoded_imm_uj[7] ),
    .B1(_19969_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _23609_ (.A0(\decoded_imm_uj[6] ),
    .A1(\mem_rdata_latched[26] ),
    .S(_19968_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _23610_ (.A0(\decoded_imm_uj[5] ),
    .A1(\mem_rdata_latched[25] ),
    .S(_19968_),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_1 _23611_ (.A0(\decoded_imm_uj[4] ),
    .A1(\mem_rdata_latched[24] ),
    .S(_19968_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _23612_ (.A0(\decoded_imm_uj[3] ),
    .A1(\mem_rdata_latched[23] ),
    .S(_19968_),
    .X(_03187_));
 sky130_fd_sc_hd__mux2_1 _23613_ (.A0(\decoded_imm_uj[2] ),
    .A1(\mem_rdata_latched[22] ),
    .S(_19968_),
    .X(_03186_));
 sky130_fd_sc_hd__buf_2 _23614_ (.A(_18577_),
    .X(_19970_));
 sky130_fd_sc_hd__mux2_1 _23615_ (.A0(\decoded_imm_uj[1] ),
    .A1(\mem_rdata_latched[21] ),
    .S(_19970_),
    .X(_03185_));
 sky130_fd_sc_hd__or3_4 _23616_ (.A(is_alu_reg_imm),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(instr_jalr),
    .X(_19971_));
 sky130_fd_sc_hd__clkbuf_2 _23617_ (.A(_19971_),
    .X(_19972_));
 sky130_fd_sc_hd__a22o_1 _23618_ (.A1(_19951_),
    .A2(\mem_rdata_q[7] ),
    .B1(_19972_),
    .B2(\mem_rdata_q[20] ),
    .X(_19973_));
 sky130_fd_sc_hd__mux2_1 _23619_ (.A0(_19973_),
    .A1(\decoded_imm[0] ),
    .S(_18905_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _23620_ (.A0(\decoded_rd[4] ),
    .A1(\mem_rdata_latched[11] ),
    .S(_19970_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _23621_ (.A0(\decoded_rd[3] ),
    .A1(\mem_rdata_latched[10] ),
    .S(_19970_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _23622_ (.A0(\decoded_rd[2] ),
    .A1(\mem_rdata_latched[9] ),
    .S(_19970_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _23623_ (.A0(\decoded_rd[1] ),
    .A1(\mem_rdata_latched[8] ),
    .S(_19970_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _23624_ (.A0(\decoded_rd[0] ),
    .A1(\mem_rdata_latched[7] ),
    .S(_19970_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_2 _23625_ (.A(instr_timer),
    .X(_19974_));
 sky130_fd_sc_hd__clkbuf_4 _23626_ (.A(_19974_),
    .X(_19975_));
 sky130_fd_sc_hd__clkbuf_2 _23627_ (.A(_18930_),
    .X(_19976_));
 sky130_fd_sc_hd__or4b_1 _23628_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[4] ),
    .D_N(\mem_rdata_q[3] ),
    .X(_19977_));
 sky130_vsdinv _23629_ (.A(\mem_rdata_q[2] ),
    .Y(_19978_));
 sky130_fd_sc_hd__and4b_2 _23630_ (.A_N(_19977_),
    .B(_19978_),
    .C(\mem_rdata_q[1] ),
    .D(\mem_rdata_q[0] ),
    .X(_19979_));
 sky130_fd_sc_hd__and3_1 _23631_ (.A(_18879_),
    .B(_18898_),
    .C(_18883_),
    .X(_19980_));
 sky130_fd_sc_hd__and3_1 _23632_ (.A(_19980_),
    .B(\mem_rdata_q[27] ),
    .C(_19954_),
    .X(_19981_));
 sky130_fd_sc_hd__a22o_1 _23633_ (.A1(_19975_),
    .A2(_19976_),
    .B1(_19979_),
    .B2(_19981_),
    .X(_03178_));
 sky130_fd_sc_hd__nor2_1 _23634_ (.A(_18589_),
    .B(_18582_),
    .Y(_19982_));
 sky130_fd_sc_hd__a22o_1 _23635_ (.A1(instr_waitirq),
    .A2(_18860_),
    .B1(_19982_),
    .B2(_19969_),
    .X(_03177_));
 sky130_vsdinv _23636_ (.A(\mem_rdata_q[28] ),
    .Y(_19983_));
 sky130_fd_sc_hd__and4_1 _23637_ (.A(_18879_),
    .B(_19983_),
    .C(\mem_rdata_q[26] ),
    .D(_18898_),
    .X(_19984_));
 sky130_fd_sc_hd__clkbuf_4 _23638_ (.A(_18713_),
    .X(_19985_));
 sky130_fd_sc_hd__a32o_1 _23639_ (.A1(_19979_),
    .A2(_18882_),
    .A3(_19984_),
    .B1(_19985_),
    .B2(_19959_),
    .X(_03176_));
 sky130_fd_sc_hd__o21ai_1 _23640_ (.A1(_18551_),
    .A2(_18578_),
    .B1(_18588_),
    .Y(_03175_));
 sky130_fd_sc_hd__a32o_1 _23641_ (.A1(_19979_),
    .A2(_19980_),
    .A3(_18882_),
    .B1(instr_setq),
    .B2(_19976_),
    .X(_03174_));
 sky130_fd_sc_hd__a22o_1 _23642_ (.A1(instr_getq),
    .A2(_19395_),
    .B1(_19979_),
    .B2(_18907_),
    .X(_03173_));
 sky130_fd_sc_hd__or4_1 _23643_ (.A(\mem_rdata_q[22] ),
    .B(\mem_rdata_q[21] ),
    .C(\mem_rdata_q[11] ),
    .D(\mem_rdata_q[10] ),
    .X(_19986_));
 sky130_fd_sc_hd__or3_1 _23644_ (.A(\mem_rdata_q[24] ),
    .B(\mem_rdata_q[23] ),
    .C(_19986_),
    .X(_19987_));
 sky130_fd_sc_hd__or4_4 _23645_ (.A(\mem_rdata_q[9] ),
    .B(\mem_rdata_q[8] ),
    .C(\mem_rdata_q[7] ),
    .D(_18927_),
    .X(_19988_));
 sky130_fd_sc_hd__nor2_2 _23646_ (.A(_19987_),
    .B(_19988_),
    .Y(_19989_));
 sky130_fd_sc_hd__or2_1 _23647_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .X(_19990_));
 sky130_fd_sc_hd__or4_4 _23648_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .D(_19990_),
    .X(_19991_));
 sky130_vsdinv _23649_ (.A(\mem_rdata_q[4] ),
    .Y(_19992_));
 sky130_fd_sc_hd__and3_1 _23650_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[1] ),
    .X(_19993_));
 sky130_fd_sc_hd__nand2_1 _23651_ (.A(_19993_),
    .B(\mem_rdata_q[0] ),
    .Y(_19994_));
 sky130_fd_sc_hd__or4_4 _23652_ (.A(_19992_),
    .B(\mem_rdata_q[3] ),
    .C(\mem_rdata_q[2] ),
    .D(_19994_),
    .X(_19995_));
 sky130_fd_sc_hd__nor2_1 _23653_ (.A(_19991_),
    .B(_19995_),
    .Y(_19996_));
 sky130_fd_sc_hd__a32o_1 _23654_ (.A1(_19989_),
    .A2(_18907_),
    .A3(_19996_),
    .B1(instr_ecall_ebreak),
    .B2(_19976_),
    .X(_03172_));
 sky130_vsdinv _23655_ (.A(\mem_rdata_q[24] ),
    .Y(_19997_));
 sky130_fd_sc_hd__and4_1 _23656_ (.A(_18878_),
    .B(_19997_),
    .C(\mem_rdata_q[31] ),
    .D(\mem_rdata_q[30] ),
    .X(_19998_));
 sky130_fd_sc_hd__nand2_1 _23657_ (.A(_19998_),
    .B(_18885_),
    .Y(_19999_));
 sky130_fd_sc_hd__or3_1 _23658_ (.A(_18919_),
    .B(_19999_),
    .C(_19991_),
    .X(_20000_));
 sky130_fd_sc_hd__or2_1 _23659_ (.A(_18880_),
    .B(_20000_),
    .X(_20001_));
 sky130_vsdinv _23660_ (.A(\mem_rdata_q[21] ),
    .Y(_20002_));
 sky130_fd_sc_hd__or4_4 _23661_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C(_18869_),
    .D(_19995_),
    .X(_20003_));
 sky130_fd_sc_hd__or3_4 _23662_ (.A(_20002_),
    .B(\mem_rdata_q[20] ),
    .C(_20003_),
    .X(_20004_));
 sky130_fd_sc_hd__buf_2 _23663_ (.A(instr_rdinstrh),
    .X(_20005_));
 sky130_fd_sc_hd__clkbuf_4 _23664_ (.A(_20005_),
    .X(_20006_));
 sky130_fd_sc_hd__buf_2 _23665_ (.A(_18908_),
    .X(_20007_));
 sky130_fd_sc_hd__a2bb2o_1 _23666_ (.A1_N(_20001_),
    .A2_N(_20004_),
    .B1(_20006_),
    .B2(_20007_),
    .X(_03171_));
 sky130_fd_sc_hd__or2_1 _23667_ (.A(\mem_rdata_q[27] ),
    .B(_20000_),
    .X(_20008_));
 sky130_fd_sc_hd__buf_2 _23668_ (.A(instr_rdinstr),
    .X(_20009_));
 sky130_fd_sc_hd__buf_2 _23669_ (.A(_20009_),
    .X(_20010_));
 sky130_fd_sc_hd__a2bb2o_1 _23670_ (.A1_N(_20008_),
    .A2_N(_20004_),
    .B1(_20010_),
    .B2(_20007_),
    .X(_03170_));
 sky130_fd_sc_hd__or2_1 _23671_ (.A(\mem_rdata_q[21] ),
    .B(_20003_),
    .X(_20011_));
 sky130_fd_sc_hd__clkbuf_4 _23672_ (.A(instr_rdcycleh),
    .X(_20012_));
 sky130_fd_sc_hd__a2bb2o_1 _23673_ (.A1_N(_20001_),
    .A2_N(_20011_),
    .B1(_20012_),
    .B2(_20007_),
    .X(_03169_));
 sky130_fd_sc_hd__a2bb2o_1 _23674_ (.A1_N(_20008_),
    .A2_N(_20011_),
    .B1(instr_rdcycle),
    .B2(_20007_),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_1 _23675_ (.A(_18932_),
    .B(_18895_),
    .Y(_20013_));
 sky130_fd_sc_hd__a22o_1 _23676_ (.A1(instr_srai),
    .A2(_19395_),
    .B1(_18901_),
    .B2(_20013_),
    .X(_03167_));
 sky130_fd_sc_hd__a22o_1 _23677_ (.A1(instr_srli),
    .A2(_19395_),
    .B1(_18907_),
    .B2(_20013_),
    .X(_03166_));
 sky130_fd_sc_hd__a32o_1 _23678_ (.A1(_18907_),
    .A2(is_alu_reg_imm),
    .A3(_18923_),
    .B1(instr_slli),
    .B2(_19976_),
    .X(_03165_));
 sky130_vsdinv _23679_ (.A(_18919_),
    .Y(_20014_));
 sky130_fd_sc_hd__and3_1 _23680_ (.A(_18881_),
    .B(_19951_),
    .C(_18592_),
    .X(_20015_));
 sky130_fd_sc_hd__a22o_1 _23681_ (.A1(instr_sw),
    .A2(_19395_),
    .B1(_20014_),
    .B2(_20015_),
    .X(_03164_));
 sky130_fd_sc_hd__a22o_1 _23682_ (.A1(_18923_),
    .A2(_20015_),
    .B1(_19959_),
    .B2(instr_sh),
    .X(_03163_));
 sky130_fd_sc_hd__a22o_1 _23683_ (.A1(_18926_),
    .A2(_20015_),
    .B1(instr_sb),
    .B2(_19976_),
    .X(_03162_));
 sky130_fd_sc_hd__and3_2 _23684_ (.A(_18881_),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(_18592_),
    .X(_20016_));
 sky130_fd_sc_hd__a22o_1 _23685_ (.A1(_18894_),
    .A2(_20016_),
    .B1(_19959_),
    .B2(instr_lhu),
    .X(_03161_));
 sky130_fd_sc_hd__a22o_1 _23686_ (.A1(_18911_),
    .A2(_20016_),
    .B1(_19959_),
    .B2(instr_lbu),
    .X(_03160_));
 sky130_fd_sc_hd__a22o_1 _23687_ (.A1(instr_lw),
    .A2(_19395_),
    .B1(_20014_),
    .B2(_20016_),
    .X(_03159_));
 sky130_fd_sc_hd__a22o_1 _23688_ (.A1(_18923_),
    .A2(_20016_),
    .B1(_19959_),
    .B2(instr_lh),
    .X(_03158_));
 sky130_fd_sc_hd__a22o_1 _23689_ (.A1(_18926_),
    .A2(_20016_),
    .B1(instr_lb),
    .B2(_19976_),
    .X(_03157_));
 sky130_fd_sc_hd__nor3_4 _23690_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .Y(_20017_));
 sky130_fd_sc_hd__and3_1 _23691_ (.A(_00325_),
    .B(_00324_),
    .C(_00326_),
    .X(_20018_));
 sky130_fd_sc_hd__and2_1 _23692_ (.A(_20018_),
    .B(_18579_),
    .X(_20019_));
 sky130_fd_sc_hd__nor2_1 _23693_ (.A(_02063_),
    .B(_18576_),
    .Y(_20020_));
 sky130_fd_sc_hd__a41o_1 _23694_ (.A1(_18578_),
    .A2(_18859_),
    .A3(_20017_),
    .A4(_20019_),
    .B1(_20020_),
    .X(_03156_));
 sky130_fd_sc_hd__nor2_1 _23695_ (.A(_00323_),
    .B(_18576_),
    .Y(_20021_));
 sky130_fd_sc_hd__a41o_1 _23696_ (.A1(_00327_),
    .A2(_18578_),
    .A3(_18859_),
    .A4(_20018_),
    .B1(_20021_),
    .X(_03155_));
 sky130_fd_sc_hd__and3_1 _23697_ (.A(_18576_),
    .B(_19940_),
    .C(_20019_),
    .X(_20022_));
 sky130_fd_sc_hd__a32o_1 _23698_ (.A1(_20022_),
    .A2(_19943_),
    .A3(_00328_),
    .B1(instr_auipc),
    .B2(_19942_),
    .X(_03154_));
 sky130_fd_sc_hd__buf_4 _23699_ (.A(instr_lui),
    .X(_20023_));
 sky130_fd_sc_hd__a32o_1 _23700_ (.A1(_20022_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(_20023_),
    .B2(_19942_),
    .X(_03153_));
 sky130_fd_sc_hd__buf_2 _23701_ (.A(\mem_rdata_q[31] ),
    .X(_20024_));
 sky130_fd_sc_hd__buf_2 _23702_ (.A(_19954_),
    .X(_20025_));
 sky130_fd_sc_hd__mux2_1 _23703_ (.A0(net298),
    .A1(_20024_),
    .S(_20025_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_1 _23704_ (.A0(net297),
    .A1(\mem_rdata_q[30] ),
    .S(_20025_),
    .X(_03151_));
 sky130_fd_sc_hd__o21a_1 _23705_ (.A1(net295),
    .A2(_19955_),
    .B1(_18897_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_4 _23706_ (.A(_19954_),
    .X(_20026_));
 sky130_fd_sc_hd__mux2_1 _23707_ (.A0(net294),
    .A1(\mem_rdata_q[28] ),
    .S(_20026_),
    .X(_03149_));
 sky130_fd_sc_hd__o21ba_1 _23708_ (.A1(net293),
    .A2(_20025_),
    .B1_N(_18882_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_1 _23709_ (.A0(net292),
    .A1(\mem_rdata_q[26] ),
    .S(_20026_),
    .X(_03147_));
 sky130_fd_sc_hd__mux2_1 _23710_ (.A0(net291),
    .A1(_18898_),
    .S(_20026_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _23711_ (.A0(net290),
    .A1(\mem_rdata_q[24] ),
    .S(_20026_),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_1 _23712_ (.A0(net289),
    .A1(\mem_rdata_q[23] ),
    .S(_20026_),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _23713_ (.A0(net288),
    .A1(\mem_rdata_q[22] ),
    .S(_20026_),
    .X(_03143_));
 sky130_fd_sc_hd__buf_4 _23714_ (.A(_19954_),
    .X(_20027_));
 sky130_fd_sc_hd__mux2_1 _23715_ (.A0(net287),
    .A1(\mem_rdata_q[21] ),
    .S(_20027_),
    .X(_03142_));
 sky130_fd_sc_hd__mux2_1 _23716_ (.A0(net286),
    .A1(\mem_rdata_q[20] ),
    .S(_20027_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_1 _23717_ (.A0(net284),
    .A1(\mem_rdata_q[19] ),
    .S(_20027_),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_1 _23718_ (.A0(net283),
    .A1(\mem_rdata_q[18] ),
    .S(_20027_),
    .X(_03139_));
 sky130_fd_sc_hd__mux2_1 _23719_ (.A0(net282),
    .A1(\mem_rdata_q[17] ),
    .S(_20027_),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_1 _23720_ (.A0(net281),
    .A1(\mem_rdata_q[16] ),
    .S(_20027_),
    .X(_03137_));
 sky130_fd_sc_hd__buf_2 _23721_ (.A(_18917_),
    .X(_20028_));
 sky130_fd_sc_hd__mux2_1 _23722_ (.A0(net280),
    .A1(\mem_rdata_q[15] ),
    .S(_20028_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_1 _23723_ (.A0(net279),
    .A1(_18893_),
    .S(_20028_),
    .X(_03135_));
 sky130_fd_sc_hd__mux2_1 _23724_ (.A0(net278),
    .A1(\mem_rdata_q[13] ),
    .S(_20028_),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_1 _23725_ (.A0(net277),
    .A1(_18889_),
    .S(_20028_),
    .X(_03133_));
 sky130_fd_sc_hd__mux2_1 _23726_ (.A0(net276),
    .A1(\mem_rdata_q[11] ),
    .S(_20028_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _23727_ (.A0(net275),
    .A1(\mem_rdata_q[10] ),
    .S(_20028_),
    .X(_03131_));
 sky130_fd_sc_hd__buf_2 _23728_ (.A(_18917_),
    .X(_20029_));
 sky130_fd_sc_hd__mux2_1 _23729_ (.A0(net305),
    .A1(\mem_rdata_q[9] ),
    .S(_20029_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_1 _23730_ (.A0(net304),
    .A1(\mem_rdata_q[8] ),
    .S(_20029_),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_1 _23731_ (.A0(net303),
    .A1(\mem_rdata_q[7] ),
    .S(_20029_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _23732_ (.A0(net302),
    .A1(\mem_rdata_q[6] ),
    .S(_20029_),
    .X(_03127_));
 sky130_fd_sc_hd__mux2_1 _23733_ (.A0(net301),
    .A1(\mem_rdata_q[5] ),
    .S(_20029_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _23734_ (.A0(net300),
    .A1(\mem_rdata_q[4] ),
    .S(_20029_),
    .X(_03125_));
 sky130_fd_sc_hd__buf_2 _23735_ (.A(_19954_),
    .X(_20030_));
 sky130_fd_sc_hd__mux2_1 _23736_ (.A0(net299),
    .A1(\mem_rdata_q[3] ),
    .S(_20030_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _23737_ (.A0(net296),
    .A1(\mem_rdata_q[2] ),
    .S(_20030_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _23738_ (.A0(net285),
    .A1(\mem_rdata_q[1] ),
    .S(_20030_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _23739_ (.A0(net274),
    .A1(\mem_rdata_q[0] ),
    .S(_20030_),
    .X(_03121_));
 sky130_vsdinv _23740_ (.A(\cpu_state[5] ),
    .Y(_20031_));
 sky130_fd_sc_hd__or3_1 _23741_ (.A(_00318_),
    .B(_00320_),
    .C(_18532_),
    .X(_20032_));
 sky130_fd_sc_hd__a31o_1 _23742_ (.A1(_18705_),
    .A2(_18722_),
    .A3(_20031_),
    .B1(_20032_),
    .X(_20033_));
 sky130_fd_sc_hd__clkbuf_4 _23743_ (.A(_20033_),
    .X(_20034_));
 sky130_fd_sc_hd__clkbuf_4 _23744_ (.A(_20034_),
    .X(_20035_));
 sky130_fd_sc_hd__mux2_1 _23745_ (.A0(_02499_),
    .A1(net330),
    .S(_20035_),
    .X(_03120_));
 sky130_fd_sc_hd__buf_4 _23746_ (.A(net329),
    .X(_20036_));
 sky130_fd_sc_hd__mux2_1 _23747_ (.A0(_02498_),
    .A1(_20036_),
    .S(_20035_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_6 _23748_ (.A(net327),
    .X(_20037_));
 sky130_fd_sc_hd__mux2_1 _23749_ (.A0(_02496_),
    .A1(_20037_),
    .S(_20035_),
    .X(_03118_));
 sky130_fd_sc_hd__buf_4 _23750_ (.A(net326),
    .X(_20038_));
 sky130_fd_sc_hd__mux2_1 _23751_ (.A0(_02495_),
    .A1(_20038_),
    .S(_20035_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _23752_ (.A0(_02494_),
    .A1(net325),
    .S(_20035_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_6 _23753_ (.A(net324),
    .X(_20039_));
 sky130_fd_sc_hd__mux2_1 _23754_ (.A0(_02493_),
    .A1(_20039_),
    .S(_20035_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_6 _23755_ (.A(net323),
    .X(_20040_));
 sky130_fd_sc_hd__buf_2 _23756_ (.A(_20034_),
    .X(_20041_));
 sky130_fd_sc_hd__mux2_1 _23757_ (.A0(_02492_),
    .A1(_20040_),
    .S(_20041_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_6 _23758_ (.A(net322),
    .X(_20042_));
 sky130_fd_sc_hd__mux2_1 _23759_ (.A0(_02491_),
    .A1(_20042_),
    .S(_20041_),
    .X(_03113_));
 sky130_fd_sc_hd__buf_6 _23760_ (.A(net321),
    .X(_20043_));
 sky130_fd_sc_hd__mux2_1 _23761_ (.A0(_02490_),
    .A1(_20043_),
    .S(_20041_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_6 _23762_ (.A(net320),
    .X(_20044_));
 sky130_fd_sc_hd__mux2_1 _23763_ (.A0(_02489_),
    .A1(_20044_),
    .S(_20041_),
    .X(_03111_));
 sky130_fd_sc_hd__buf_6 _23764_ (.A(net319),
    .X(_20045_));
 sky130_fd_sc_hd__mux2_1 _23765_ (.A0(_02488_),
    .A1(_20045_),
    .S(_20041_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_6 _23766_ (.A(net318),
    .X(_20046_));
 sky130_fd_sc_hd__mux2_1 _23767_ (.A0(_02487_),
    .A1(_20046_),
    .S(_20041_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_6 _23768_ (.A(net316),
    .X(_20047_));
 sky130_fd_sc_hd__clkbuf_4 _23769_ (.A(_20034_),
    .X(_20048_));
 sky130_fd_sc_hd__mux2_1 _23770_ (.A0(_02485_),
    .A1(_20047_),
    .S(_20048_),
    .X(_03108_));
 sky130_fd_sc_hd__buf_6 _23771_ (.A(net315),
    .X(_20049_));
 sky130_fd_sc_hd__mux2_1 _23772_ (.A0(_02484_),
    .A1(_20049_),
    .S(_20048_),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _23773_ (.A0(_02483_),
    .A1(net314),
    .S(_20048_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_4 _23774_ (.A(net313),
    .X(_20050_));
 sky130_fd_sc_hd__mux2_1 _23775_ (.A0(_02482_),
    .A1(_20050_),
    .S(_20048_),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _23776_ (.A0(_02481_),
    .A1(net312),
    .S(_20048_),
    .X(_03104_));
 sky130_fd_sc_hd__buf_4 _23777_ (.A(net311),
    .X(_20051_));
 sky130_fd_sc_hd__mux2_1 _23778_ (.A0(_02480_),
    .A1(_20051_),
    .S(_20048_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_2 _23779_ (.A(_20034_),
    .X(_20052_));
 sky130_fd_sc_hd__mux2_1 _23780_ (.A0(_02479_),
    .A1(net310),
    .S(_20052_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_2 _23781_ (.A(net309),
    .X(_20053_));
 sky130_fd_sc_hd__mux2_1 _23782_ (.A0(_02478_),
    .A1(_20053_),
    .S(_20052_),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _23783_ (.A0(_02477_),
    .A1(net308),
    .S(_20052_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_4 _23784_ (.A(net307),
    .X(_20054_));
 sky130_fd_sc_hd__mux2_1 _23785_ (.A0(_02476_),
    .A1(_20054_),
    .S(_20052_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_2 _23786_ (.A(net337),
    .X(_20055_));
 sky130_fd_sc_hd__mux2_1 _23787_ (.A0(_02506_),
    .A1(_20055_),
    .S(_20052_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_2 _23788_ (.A(net336),
    .X(_20056_));
 sky130_fd_sc_hd__mux2_1 _23789_ (.A0(_02505_),
    .A1(_20056_),
    .S(_20052_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_4 _23790_ (.A(net335),
    .X(_20057_));
 sky130_fd_sc_hd__buf_2 _23791_ (.A(_20033_),
    .X(_20058_));
 sky130_fd_sc_hd__mux2_1 _23792_ (.A0(_02504_),
    .A1(_20057_),
    .S(_20058_),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_1 _23793_ (.A0(_02503_),
    .A1(net334),
    .S(_20058_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_4 _23794_ (.A(net333),
    .X(_20059_));
 sky130_fd_sc_hd__mux2_1 _23795_ (.A0(_02502_),
    .A1(_20059_),
    .S(_20058_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_4 _23796_ (.A(net332),
    .X(_20060_));
 sky130_fd_sc_hd__mux2_1 _23797_ (.A0(_02501_),
    .A1(_20060_),
    .S(_20058_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_4 _23798_ (.A(net331),
    .X(_20061_));
 sky130_fd_sc_hd__mux2_1 _23799_ (.A0(_02500_),
    .A1(_20061_),
    .S(_20058_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_4 _23800_ (.A(net328),
    .X(_20062_));
 sky130_fd_sc_hd__mux2_1 _23801_ (.A0(_02497_),
    .A1(_20062_),
    .S(_20058_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_8 _23802_ (.A(net317),
    .X(_20063_));
 sky130_fd_sc_hd__mux2_1 _23803_ (.A0(_02486_),
    .A1(_20063_),
    .S(_20034_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_6 _23804_ (.A(net306),
    .X(_20064_));
 sky130_fd_sc_hd__mux2_1 _23805_ (.A0(_02475_),
    .A1(_20064_),
    .S(_20034_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _23806_ (.A0(net158),
    .A1(net191),
    .S(net425),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _23807_ (.A0(net157),
    .A1(net190),
    .S(_18857_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _23808_ (.A0(net155),
    .A1(net188),
    .S(net425),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _23809_ (.A0(net154),
    .A1(net187),
    .S(net425),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_1 _23810_ (.A0(net153),
    .A1(net186),
    .S(_18857_),
    .X(_03084_));
 sky130_fd_sc_hd__buf_2 _23811_ (.A(net427),
    .X(_20065_));
 sky130_fd_sc_hd__mux2_1 _23812_ (.A0(net152),
    .A1(net185),
    .S(net420),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _23813_ (.A0(net151),
    .A1(net184),
    .S(net420),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _23814_ (.A0(net150),
    .A1(net183),
    .S(net420),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _23815_ (.A0(net149),
    .A1(net182),
    .S(net420),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_1 _23816_ (.A0(net148),
    .A1(net181),
    .S(_20065_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _23817_ (.A0(net147),
    .A1(net180),
    .S(net420),
    .X(_03078_));
 sky130_fd_sc_hd__buf_6 _23818_ (.A(net427),
    .X(_20066_));
 sky130_fd_sc_hd__mux2_1 _23819_ (.A0(net146),
    .A1(net179),
    .S(net419),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _23820_ (.A0(net144),
    .A1(net177),
    .S(net419),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _23821_ (.A0(net143),
    .A1(net176),
    .S(net419),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_1 _23822_ (.A0(net142),
    .A1(net175),
    .S(_20066_),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_1 _23823_ (.A0(net141),
    .A1(net174),
    .S(_20066_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _23824_ (.A0(net140),
    .A1(net173),
    .S(net419),
    .X(_03072_));
 sky130_fd_sc_hd__buf_1 _23825_ (.A(net427),
    .X(_20067_));
 sky130_fd_sc_hd__mux2_1 _23826_ (.A0(net139),
    .A1(net172),
    .S(net418),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _23827_ (.A0(net138),
    .A1(net171),
    .S(net417),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _23828_ (.A0(net137),
    .A1(net170),
    .S(net417),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_1 _23829_ (.A0(net136),
    .A1(net169),
    .S(net417),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _23830_ (.A0(net135),
    .A1(net168),
    .S(_20067_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_1 _23831_ (.A0(net165),
    .A1(net198),
    .S(net418),
    .X(_03066_));
 sky130_fd_sc_hd__buf_2 _23832_ (.A(_18856_),
    .X(_20068_));
 sky130_fd_sc_hd__mux2_1 _23833_ (.A0(net164),
    .A1(net197),
    .S(net416),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _23834_ (.A0(net163),
    .A1(net196),
    .S(net416),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_1 _23835_ (.A0(net162),
    .A1(net195),
    .S(net416),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _23836_ (.A0(net161),
    .A1(net194),
    .S(net416),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _23837_ (.A0(net160),
    .A1(net193),
    .S(net416),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _23838_ (.A0(net159),
    .A1(net192),
    .S(net416),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _23839_ (.A0(net156),
    .A1(net189),
    .S(net427),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_4 _23840_ (.A(\pcpi_mul.rs1[31] ),
    .X(_20069_));
 sky130_fd_sc_hd__buf_6 _23841_ (.A(_20069_),
    .X(_20070_));
 sky130_fd_sc_hd__buf_6 _23842_ (.A(_20070_),
    .X(_20071_));
 sky130_fd_sc_hd__a21o_1 _23843_ (.A1(_20071_),
    .A2(_18689_),
    .B1(_18681_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_6 _23844_ (.A(\pcpi_mul.rs1[30] ),
    .X(_20072_));
 sky130_fd_sc_hd__clkbuf_4 _23845_ (.A(_20072_),
    .X(_20073_));
 sky130_fd_sc_hd__buf_4 _23846_ (.A(_20073_),
    .X(_20074_));
 sky130_fd_sc_hd__buf_2 _23847_ (.A(_20074_),
    .X(_20075_));
 sky130_fd_sc_hd__buf_2 _23848_ (.A(_19883_),
    .X(_20076_));
 sky130_fd_sc_hd__mux2_1 _23849_ (.A0(_20036_),
    .A1(_20075_),
    .S(_20076_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_4 _23850_ (.A(\pcpi_mul.rs1[29] ),
    .X(_20077_));
 sky130_fd_sc_hd__buf_4 _23851_ (.A(_20077_),
    .X(_20078_));
 sky130_fd_sc_hd__buf_4 _23852_ (.A(_20078_),
    .X(_20079_));
 sky130_fd_sc_hd__buf_2 _23853_ (.A(_20079_),
    .X(_20080_));
 sky130_fd_sc_hd__mux2_1 _23854_ (.A0(_20037_),
    .A1(_20080_),
    .S(_20076_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_4 _23855_ (.A(\pcpi_mul.rs1[28] ),
    .X(_20081_));
 sky130_fd_sc_hd__buf_6 _23856_ (.A(_20081_),
    .X(_20082_));
 sky130_fd_sc_hd__clkbuf_4 _23857_ (.A(_20082_),
    .X(_20083_));
 sky130_fd_sc_hd__clkbuf_4 _23858_ (.A(_20083_),
    .X(_20084_));
 sky130_fd_sc_hd__mux2_1 _23859_ (.A0(_20038_),
    .A1(_20084_),
    .S(_20076_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_2 _23860_ (.A(\pcpi_mul.rs1[27] ),
    .X(_20085_));
 sky130_fd_sc_hd__buf_4 _23861_ (.A(_20085_),
    .X(_20086_));
 sky130_fd_sc_hd__buf_6 _23862_ (.A(_20086_),
    .X(_20087_));
 sky130_fd_sc_hd__clkbuf_4 _23863_ (.A(_20087_),
    .X(_20088_));
 sky130_fd_sc_hd__clkbuf_4 _23864_ (.A(_20088_),
    .X(_20089_));
 sky130_fd_sc_hd__mux2_1 _23865_ (.A0(net325),
    .A1(_20089_),
    .S(_20076_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_4 _23866_ (.A(\pcpi_mul.rs1[26] ),
    .X(_20090_));
 sky130_fd_sc_hd__buf_4 _23867_ (.A(_20090_),
    .X(_20091_));
 sky130_fd_sc_hd__clkbuf_4 _23868_ (.A(_20091_),
    .X(_20092_));
 sky130_fd_sc_hd__mux2_1 _23869_ (.A0(_20039_),
    .A1(_20092_),
    .S(_20076_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_4 _23870_ (.A(\pcpi_mul.rs1[25] ),
    .X(_20093_));
 sky130_fd_sc_hd__buf_4 _23871_ (.A(_20093_),
    .X(_20094_));
 sky130_fd_sc_hd__clkbuf_4 _23872_ (.A(_20094_),
    .X(_20095_));
 sky130_fd_sc_hd__mux2_1 _23873_ (.A0(_20040_),
    .A1(_20095_),
    .S(_20076_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_2 _23874_ (.A(\pcpi_mul.rs1[24] ),
    .X(_20096_));
 sky130_fd_sc_hd__clkbuf_4 _23875_ (.A(_20096_),
    .X(_20097_));
 sky130_fd_sc_hd__buf_4 _23876_ (.A(_20097_),
    .X(_20098_));
 sky130_fd_sc_hd__buf_2 _23877_ (.A(_20098_),
    .X(_20099_));
 sky130_fd_sc_hd__buf_2 _23878_ (.A(_19883_),
    .X(_20100_));
 sky130_fd_sc_hd__mux2_1 _23879_ (.A0(_20042_),
    .A1(_20099_),
    .S(_20100_),
    .X(_03051_));
 sky130_fd_sc_hd__buf_4 _23880_ (.A(\pcpi_mul.rs1[23] ),
    .X(_20101_));
 sky130_fd_sc_hd__buf_4 _23881_ (.A(_20101_),
    .X(_20102_));
 sky130_fd_sc_hd__buf_4 _23882_ (.A(_20102_),
    .X(_20103_));
 sky130_fd_sc_hd__mux2_1 _23883_ (.A0(_20043_),
    .A1(_20103_),
    .S(_20100_),
    .X(_03050_));
 sky130_fd_sc_hd__buf_4 _23884_ (.A(\pcpi_mul.rs1[22] ),
    .X(_20104_));
 sky130_fd_sc_hd__buf_4 _23885_ (.A(_20104_),
    .X(_20105_));
 sky130_fd_sc_hd__buf_2 _23886_ (.A(_20105_),
    .X(_20106_));
 sky130_fd_sc_hd__mux2_1 _23887_ (.A0(_20044_),
    .A1(_20106_),
    .S(_20100_),
    .X(_03049_));
 sky130_fd_sc_hd__buf_6 _23888_ (.A(\pcpi_mul.rs1[21] ),
    .X(_20107_));
 sky130_fd_sc_hd__buf_6 _23889_ (.A(_20107_),
    .X(_20108_));
 sky130_fd_sc_hd__buf_2 _23890_ (.A(_20108_),
    .X(_20109_));
 sky130_fd_sc_hd__mux2_1 _23891_ (.A0(_20045_),
    .A1(_20109_),
    .S(_20100_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_4 _23892_ (.A(\pcpi_mul.rs1[20] ),
    .X(_20110_));
 sky130_fd_sc_hd__buf_4 _23893_ (.A(_20110_),
    .X(_20111_));
 sky130_fd_sc_hd__clkbuf_4 _23894_ (.A(_20111_),
    .X(_20112_));
 sky130_fd_sc_hd__mux2_1 _23895_ (.A0(_20046_),
    .A1(_20112_),
    .S(_20100_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_4 _23896_ (.A(\pcpi_mul.rs1[19] ),
    .X(_20113_));
 sky130_fd_sc_hd__buf_4 _23897_ (.A(_20113_),
    .X(_20114_));
 sky130_fd_sc_hd__buf_4 _23898_ (.A(_20114_),
    .X(_20115_));
 sky130_fd_sc_hd__buf_4 _23899_ (.A(_20115_),
    .X(_20116_));
 sky130_fd_sc_hd__mux2_1 _23900_ (.A0(_20047_),
    .A1(_20116_),
    .S(_20100_),
    .X(_03046_));
 sky130_fd_sc_hd__buf_2 _23901_ (.A(\pcpi_mul.rs1[18] ),
    .X(_20117_));
 sky130_fd_sc_hd__clkbuf_4 _23902_ (.A(_20117_),
    .X(_20118_));
 sky130_fd_sc_hd__clkbuf_4 _23903_ (.A(_20118_),
    .X(_20119_));
 sky130_fd_sc_hd__buf_4 _23904_ (.A(_20119_),
    .X(_20120_));
 sky130_fd_sc_hd__buf_2 _23905_ (.A(_19883_),
    .X(_20121_));
 sky130_fd_sc_hd__mux2_1 _23906_ (.A0(_20049_),
    .A1(_20120_),
    .S(_20121_),
    .X(_03045_));
 sky130_fd_sc_hd__buf_4 _23907_ (.A(\pcpi_mul.rs1[17] ),
    .X(_20122_));
 sky130_fd_sc_hd__clkbuf_4 _23908_ (.A(_20122_),
    .X(_20123_));
 sky130_fd_sc_hd__buf_4 _23909_ (.A(_20123_),
    .X(_20124_));
 sky130_fd_sc_hd__mux2_1 _23910_ (.A0(net314),
    .A1(_20124_),
    .S(_20121_),
    .X(_03044_));
 sky130_fd_sc_hd__buf_4 _23911_ (.A(\pcpi_mul.rs1[16] ),
    .X(_20125_));
 sky130_fd_sc_hd__buf_6 _23912_ (.A(_20125_),
    .X(_20126_));
 sky130_fd_sc_hd__clkbuf_8 _23913_ (.A(_20126_),
    .X(_20127_));
 sky130_fd_sc_hd__mux2_1 _23914_ (.A0(_20050_),
    .A1(_20127_),
    .S(_20121_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_4 _23915_ (.A(\pcpi_mul.rs1[15] ),
    .X(_20128_));
 sky130_fd_sc_hd__buf_4 _23916_ (.A(_20128_),
    .X(_20129_));
 sky130_fd_sc_hd__buf_6 _23917_ (.A(_20129_),
    .X(_20130_));
 sky130_fd_sc_hd__buf_8 _23918_ (.A(_20130_),
    .X(_20131_));
 sky130_fd_sc_hd__mux2_1 _23919_ (.A0(net312),
    .A1(_20131_),
    .S(_20121_),
    .X(_03042_));
 sky130_fd_sc_hd__buf_6 _23920_ (.A(\pcpi_mul.rs1[14] ),
    .X(_20132_));
 sky130_fd_sc_hd__buf_4 _23921_ (.A(_20132_),
    .X(_20133_));
 sky130_fd_sc_hd__buf_8 _23922_ (.A(_20133_),
    .X(_20134_));
 sky130_fd_sc_hd__mux2_1 _23923_ (.A0(_20051_),
    .A1(_20134_),
    .S(_20121_),
    .X(_03041_));
 sky130_fd_sc_hd__buf_4 _23924_ (.A(\pcpi_mul.rs1[13] ),
    .X(_20135_));
 sky130_fd_sc_hd__buf_6 _23925_ (.A(_20135_),
    .X(_20136_));
 sky130_fd_sc_hd__mux2_1 _23926_ (.A0(net310),
    .A1(_20136_),
    .S(_20121_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_4 _23927_ (.A(\pcpi_mul.rs1[12] ),
    .X(_20137_));
 sky130_fd_sc_hd__buf_8 _23928_ (.A(_20137_),
    .X(_20138_));
 sky130_fd_sc_hd__clkbuf_8 _23929_ (.A(_20138_),
    .X(_20139_));
 sky130_fd_sc_hd__buf_2 _23930_ (.A(_18679_),
    .X(_20140_));
 sky130_fd_sc_hd__mux2_1 _23931_ (.A0(_20053_),
    .A1(_20139_),
    .S(_20140_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_4 _23932_ (.A(\pcpi_mul.rs1[11] ),
    .X(_20141_));
 sky130_fd_sc_hd__buf_6 _23933_ (.A(_20141_),
    .X(_20142_));
 sky130_fd_sc_hd__clkbuf_8 _23934_ (.A(_20142_),
    .X(_20143_));
 sky130_fd_sc_hd__mux2_1 _23935_ (.A0(net308),
    .A1(_20143_),
    .S(_20140_),
    .X(_03038_));
 sky130_fd_sc_hd__buf_4 _23936_ (.A(\pcpi_mul.rs1[10] ),
    .X(_20144_));
 sky130_fd_sc_hd__buf_6 _23937_ (.A(_20144_),
    .X(_20145_));
 sky130_fd_sc_hd__buf_6 _23938_ (.A(_20145_),
    .X(_20146_));
 sky130_fd_sc_hd__buf_8 _23939_ (.A(_20146_),
    .X(_20147_));
 sky130_fd_sc_hd__mux2_1 _23940_ (.A0(_20054_),
    .A1(_20147_),
    .S(_20140_),
    .X(_03037_));
 sky130_fd_sc_hd__buf_8 _23941_ (.A(\pcpi_mul.rs1[9] ),
    .X(_20148_));
 sky130_fd_sc_hd__buf_4 _23942_ (.A(_20148_),
    .X(_20149_));
 sky130_fd_sc_hd__buf_1 _23943_ (.A(_20149_),
    .X(_20150_));
 sky130_fd_sc_hd__mux2_1 _23944_ (.A0(_20055_),
    .A1(net454),
    .S(_20140_),
    .X(_03036_));
 sky130_fd_sc_hd__buf_6 _23945_ (.A(\pcpi_mul.rs1[8] ),
    .X(_20151_));
 sky130_fd_sc_hd__buf_6 _23946_ (.A(_20151_),
    .X(_20152_));
 sky130_fd_sc_hd__clkbuf_8 _23947_ (.A(_20152_),
    .X(_20153_));
 sky130_fd_sc_hd__mux2_1 _23948_ (.A0(_20056_),
    .A1(_20153_),
    .S(_20140_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_4 _23949_ (.A(\pcpi_mul.rs1[7] ),
    .X(_20154_));
 sky130_fd_sc_hd__buf_4 _23950_ (.A(_20154_),
    .X(_20155_));
 sky130_fd_sc_hd__buf_6 _23951_ (.A(_20155_),
    .X(_20156_));
 sky130_fd_sc_hd__buf_6 _23952_ (.A(_20156_),
    .X(_20157_));
 sky130_fd_sc_hd__mux2_1 _23953_ (.A0(_20057_),
    .A1(_20157_),
    .S(_20140_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_4 _23954_ (.A(\pcpi_mul.rs1[6] ),
    .X(_20158_));
 sky130_fd_sc_hd__buf_6 _23955_ (.A(_20158_),
    .X(_20159_));
 sky130_fd_sc_hd__clkbuf_4 _23956_ (.A(_18679_),
    .X(_20160_));
 sky130_fd_sc_hd__mux2_1 _23957_ (.A0(net334),
    .A1(_20159_),
    .S(_20160_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_4 _23958_ (.A(\pcpi_mul.rs1[5] ),
    .X(_20161_));
 sky130_fd_sc_hd__buf_6 _23959_ (.A(_20161_),
    .X(_20162_));
 sky130_fd_sc_hd__buf_6 _23960_ (.A(_20162_),
    .X(_20163_));
 sky130_fd_sc_hd__mux2_1 _23961_ (.A0(_20059_),
    .A1(_20163_),
    .S(_20160_),
    .X(_03032_));
 sky130_fd_sc_hd__buf_4 _23962_ (.A(\pcpi_mul.rs1[4] ),
    .X(_20164_));
 sky130_fd_sc_hd__buf_4 _23963_ (.A(_20164_),
    .X(_20165_));
 sky130_fd_sc_hd__buf_6 _23964_ (.A(_20165_),
    .X(_20166_));
 sky130_fd_sc_hd__mux2_1 _23965_ (.A0(_20060_),
    .A1(_20166_),
    .S(_20160_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_4 _23966_ (.A(\pcpi_mul.rs1[3] ),
    .X(_20167_));
 sky130_fd_sc_hd__buf_6 _23967_ (.A(_20167_),
    .X(_20168_));
 sky130_fd_sc_hd__buf_6 _23968_ (.A(_20168_),
    .X(_20169_));
 sky130_fd_sc_hd__mux2_1 _23969_ (.A0(_20061_),
    .A1(_20169_),
    .S(_20160_),
    .X(_03030_));
 sky130_fd_sc_hd__buf_6 _23970_ (.A(\pcpi_mul.rs1[2] ),
    .X(_20170_));
 sky130_fd_sc_hd__buf_6 _23971_ (.A(_20170_),
    .X(_20171_));
 sky130_fd_sc_hd__buf_6 _23972_ (.A(_20171_),
    .X(_20172_));
 sky130_fd_sc_hd__mux2_1 _23973_ (.A0(_20062_),
    .A1(_20172_),
    .S(_20160_),
    .X(_03029_));
 sky130_fd_sc_hd__buf_4 _23974_ (.A(\pcpi_mul.rs1[1] ),
    .X(_20173_));
 sky130_fd_sc_hd__clkbuf_4 _23975_ (.A(_20173_),
    .X(_20174_));
 sky130_fd_sc_hd__buf_4 _23976_ (.A(_20174_),
    .X(_20175_));
 sky130_fd_sc_hd__mux2_1 _23977_ (.A0(_20063_),
    .A1(_20175_),
    .S(_20160_),
    .X(_03028_));
 sky130_fd_sc_hd__buf_4 _23978_ (.A(\pcpi_mul.rs1[0] ),
    .X(_20176_));
 sky130_fd_sc_hd__buf_6 _23979_ (.A(_20176_),
    .X(_20177_));
 sky130_fd_sc_hd__buf_6 _23980_ (.A(_20177_),
    .X(_20178_));
 sky130_fd_sc_hd__mux2_1 _23981_ (.A0(_20064_),
    .A1(_20178_),
    .S(_18680_),
    .X(_03027_));
 sky130_fd_sc_hd__nand2_1 _23982_ (.A(_19642_),
    .B(_19603_),
    .Y(_20179_));
 sky130_fd_sc_hd__buf_6 _23983_ (.A(_20179_),
    .X(_20180_));
 sky130_fd_sc_hd__buf_4 _23984_ (.A(_20180_),
    .X(_20181_));
 sky130_fd_sc_hd__mux2_1 _23985_ (.A0(_19720_),
    .A1(\cpuregs[5][31] ),
    .S(_20181_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _23986_ (.A0(_19724_),
    .A1(\cpuregs[5][30] ),
    .S(_20181_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_1 _23987_ (.A0(_19725_),
    .A1(\cpuregs[5][29] ),
    .S(_20181_),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_1 _23988_ (.A0(_19726_),
    .A1(\cpuregs[5][28] ),
    .S(_20181_),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_1 _23989_ (.A0(_19727_),
    .A1(\cpuregs[5][27] ),
    .S(_20181_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _23990_ (.A0(_19728_),
    .A1(\cpuregs[5][26] ),
    .S(_20181_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_4 _23991_ (.A(_20180_),
    .X(_20182_));
 sky130_fd_sc_hd__mux2_1 _23992_ (.A0(_19729_),
    .A1(\cpuregs[5][25] ),
    .S(_20182_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _23993_ (.A0(_19731_),
    .A1(\cpuregs[5][24] ),
    .S(_20182_),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_1 _23994_ (.A0(_19732_),
    .A1(\cpuregs[5][23] ),
    .S(_20182_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _23995_ (.A0(_19733_),
    .A1(\cpuregs[5][22] ),
    .S(_20182_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _23996_ (.A0(_19734_),
    .A1(\cpuregs[5][21] ),
    .S(_20182_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _23997_ (.A0(_19735_),
    .A1(\cpuregs[5][20] ),
    .S(_20182_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_4 _23998_ (.A(_20180_),
    .X(_20183_));
 sky130_fd_sc_hd__mux2_1 _23999_ (.A0(_19736_),
    .A1(\cpuregs[5][19] ),
    .S(_20183_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _24000_ (.A0(_19738_),
    .A1(\cpuregs[5][18] ),
    .S(_20183_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _24001_ (.A0(_19739_),
    .A1(\cpuregs[5][17] ),
    .S(_20183_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _24002_ (.A0(_19740_),
    .A1(\cpuregs[5][16] ),
    .S(_20183_),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_1 _24003_ (.A0(_19741_),
    .A1(\cpuregs[5][15] ),
    .S(_20183_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _24004_ (.A0(_19742_),
    .A1(\cpuregs[5][14] ),
    .S(_20183_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_4 _24005_ (.A(_20180_),
    .X(_20184_));
 sky130_fd_sc_hd__mux2_1 _24006_ (.A0(_19743_),
    .A1(\cpuregs[5][13] ),
    .S(_20184_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _24007_ (.A0(_19745_),
    .A1(\cpuregs[5][12] ),
    .S(_20184_),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _24008_ (.A0(_19746_),
    .A1(\cpuregs[5][11] ),
    .S(_20184_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _24009_ (.A0(_19747_),
    .A1(\cpuregs[5][10] ),
    .S(_20184_),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_1 _24010_ (.A0(_19748_),
    .A1(\cpuregs[5][9] ),
    .S(_20184_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _24011_ (.A0(_19749_),
    .A1(\cpuregs[5][8] ),
    .S(_20184_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_4 _24012_ (.A(_20179_),
    .X(_20185_));
 sky130_fd_sc_hd__mux2_1 _24013_ (.A0(_19750_),
    .A1(\cpuregs[5][7] ),
    .S(_20185_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_1 _24014_ (.A0(_19752_),
    .A1(\cpuregs[5][6] ),
    .S(_20185_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_1 _24015_ (.A0(_19753_),
    .A1(\cpuregs[5][5] ),
    .S(_20185_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _24016_ (.A0(_19754_),
    .A1(\cpuregs[5][4] ),
    .S(_20185_),
    .X(_02999_));
 sky130_fd_sc_hd__mux2_1 _24017_ (.A0(_19755_),
    .A1(\cpuregs[5][3] ),
    .S(_20185_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_1 _24018_ (.A0(_19756_),
    .A1(\cpuregs[5][2] ),
    .S(_20185_),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_1 _24019_ (.A0(_19757_),
    .A1(\cpuregs[5][1] ),
    .S(_20180_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _24020_ (.A0(_19758_),
    .A1(\cpuregs[5][0] ),
    .S(_20180_),
    .X(_02995_));
 sky130_fd_sc_hd__nand2_1 _24021_ (.A(_19601_),
    .B(_19759_),
    .Y(_20186_));
 sky130_fd_sc_hd__buf_6 _24022_ (.A(_20186_),
    .X(_20187_));
 sky130_fd_sc_hd__buf_4 _24023_ (.A(_20187_),
    .X(_20188_));
 sky130_fd_sc_hd__mux2_1 _24024_ (.A0(_19720_),
    .A1(\cpuregs[2][31] ),
    .S(_20188_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _24025_ (.A0(_19724_),
    .A1(\cpuregs[2][30] ),
    .S(_20188_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _24026_ (.A0(_19725_),
    .A1(\cpuregs[2][29] ),
    .S(_20188_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _24027_ (.A0(_19726_),
    .A1(\cpuregs[2][28] ),
    .S(_20188_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _24028_ (.A0(_19727_),
    .A1(\cpuregs[2][27] ),
    .S(_20188_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _24029_ (.A0(_19728_),
    .A1(\cpuregs[2][26] ),
    .S(_20188_),
    .X(_02989_));
 sky130_fd_sc_hd__buf_4 _24030_ (.A(_20187_),
    .X(_20189_));
 sky130_fd_sc_hd__mux2_1 _24031_ (.A0(_19729_),
    .A1(\cpuregs[2][25] ),
    .S(_20189_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _24032_ (.A0(_19731_),
    .A1(\cpuregs[2][24] ),
    .S(_20189_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _24033_ (.A0(_19732_),
    .A1(\cpuregs[2][23] ),
    .S(_20189_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _24034_ (.A0(_19733_),
    .A1(\cpuregs[2][22] ),
    .S(_20189_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _24035_ (.A0(_19734_),
    .A1(\cpuregs[2][21] ),
    .S(_20189_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _24036_ (.A0(_19735_),
    .A1(\cpuregs[2][20] ),
    .S(_20189_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_4 _24037_ (.A(_20187_),
    .X(_20190_));
 sky130_fd_sc_hd__mux2_1 _24038_ (.A0(_19736_),
    .A1(\cpuregs[2][19] ),
    .S(_20190_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _24039_ (.A0(_19738_),
    .A1(\cpuregs[2][18] ),
    .S(_20190_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _24040_ (.A0(_19739_),
    .A1(\cpuregs[2][17] ),
    .S(_20190_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _24041_ (.A0(_19740_),
    .A1(\cpuregs[2][16] ),
    .S(_20190_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _24042_ (.A0(_19741_),
    .A1(\cpuregs[2][15] ),
    .S(_20190_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _24043_ (.A0(_19742_),
    .A1(\cpuregs[2][14] ),
    .S(_20190_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_4 _24044_ (.A(_20187_),
    .X(_20191_));
 sky130_fd_sc_hd__mux2_1 _24045_ (.A0(_19743_),
    .A1(\cpuregs[2][13] ),
    .S(_20191_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _24046_ (.A0(_19745_),
    .A1(\cpuregs[2][12] ),
    .S(_20191_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _24047_ (.A0(_19746_),
    .A1(\cpuregs[2][11] ),
    .S(_20191_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _24048_ (.A0(_19747_),
    .A1(\cpuregs[2][10] ),
    .S(_20191_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _24049_ (.A0(_19748_),
    .A1(\cpuregs[2][9] ),
    .S(_20191_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _24050_ (.A0(_19749_),
    .A1(\cpuregs[2][8] ),
    .S(_20191_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_4 _24051_ (.A(_20186_),
    .X(_20192_));
 sky130_fd_sc_hd__mux2_1 _24052_ (.A0(_19750_),
    .A1(\cpuregs[2][7] ),
    .S(_20192_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _24053_ (.A0(_19752_),
    .A1(\cpuregs[2][6] ),
    .S(_20192_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _24054_ (.A0(_19753_),
    .A1(\cpuregs[2][5] ),
    .S(_20192_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _24055_ (.A0(_19754_),
    .A1(\cpuregs[2][4] ),
    .S(_20192_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _24056_ (.A0(_19755_),
    .A1(\cpuregs[2][3] ),
    .S(_20192_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _24057_ (.A0(_19756_),
    .A1(\cpuregs[2][2] ),
    .S(_20192_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _24058_ (.A0(_19757_),
    .A1(\cpuregs[2][1] ),
    .S(_20187_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _24059_ (.A0(_19758_),
    .A1(\cpuregs[2][0] ),
    .S(_20187_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_4 _24060_ (.A(_18527_),
    .X(_20193_));
 sky130_vsdinv _24061_ (.A(_20193_),
    .Y(mem_xfer));
 sky130_fd_sc_hd__mux2_1 _24062_ (.A0(net57),
    .A1(_20024_),
    .S(_20193_),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _24063_ (.A0(net523),
    .A1(\mem_rdata_q[30] ),
    .S(_20193_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _24064_ (.A0(net54),
    .A1(\mem_rdata_q[29] ),
    .S(_20193_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _24065_ (.A0(net53),
    .A1(\mem_rdata_q[28] ),
    .S(_20193_),
    .X(_02959_));
 sky130_fd_sc_hd__buf_2 _24066_ (.A(_18527_),
    .X(_20194_));
 sky130_fd_sc_hd__clkbuf_4 _24067_ (.A(_20194_),
    .X(_20195_));
 sky130_fd_sc_hd__mux2_1 _24068_ (.A0(net52),
    .A1(\mem_rdata_q[27] ),
    .S(_20195_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _24069_ (.A0(net51),
    .A1(\mem_rdata_q[26] ),
    .S(_20195_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _24070_ (.A0(net50),
    .A1(_18898_),
    .S(_20195_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _24071_ (.A0(net49),
    .A1(\mem_rdata_q[24] ),
    .S(_20195_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_1 _24072_ (.A0(net48),
    .A1(\mem_rdata_q[23] ),
    .S(_20195_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _24073_ (.A0(net47),
    .A1(\mem_rdata_q[22] ),
    .S(_20195_),
    .X(_02953_));
 sky130_fd_sc_hd__buf_2 _24074_ (.A(_20194_),
    .X(_20196_));
 sky130_fd_sc_hd__mux2_1 _24075_ (.A0(net46),
    .A1(\mem_rdata_q[21] ),
    .S(_20196_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _24076_ (.A0(net524),
    .A1(\mem_rdata_q[20] ),
    .S(_20196_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _24077_ (.A0(net526),
    .A1(\mem_rdata_q[19] ),
    .S(_20196_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _24078_ (.A0(net42),
    .A1(\mem_rdata_q[18] ),
    .S(_20196_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _24079_ (.A0(net41),
    .A1(\mem_rdata_q[17] ),
    .S(_20196_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _24080_ (.A0(net40),
    .A1(\mem_rdata_q[16] ),
    .S(_20196_),
    .X(_02947_));
 sky130_fd_sc_hd__buf_2 _24081_ (.A(_18527_),
    .X(_20197_));
 sky130_fd_sc_hd__mux2_1 _24082_ (.A0(net527),
    .A1(\mem_rdata_q[15] ),
    .S(_20197_),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_1 _24083_ (.A0(net38),
    .A1(_18893_),
    .S(_20197_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _24084_ (.A0(net37),
    .A1(\mem_rdata_q[13] ),
    .S(_20197_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _24085_ (.A0(net528),
    .A1(_18889_),
    .S(_20197_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _24086_ (.A0(net35),
    .A1(\mem_rdata_q[11] ),
    .S(_20197_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _24087_ (.A0(net34),
    .A1(\mem_rdata_q[10] ),
    .S(_20197_),
    .X(_02941_));
 sky130_fd_sc_hd__buf_2 _24088_ (.A(_18527_),
    .X(_20198_));
 sky130_fd_sc_hd__mux2_1 _24089_ (.A0(net64),
    .A1(\mem_rdata_q[9] ),
    .S(_20198_),
    .X(_02940_));
 sky130_fd_sc_hd__mux2_1 _24090_ (.A0(net63),
    .A1(\mem_rdata_q[8] ),
    .S(_20198_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _24091_ (.A0(net62),
    .A1(\mem_rdata_q[7] ),
    .S(_20198_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _24092_ (.A0(net61),
    .A1(\mem_rdata_q[6] ),
    .S(_20198_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _24093_ (.A0(net522),
    .A1(\mem_rdata_q[5] ),
    .S(_20198_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _24094_ (.A0(net59),
    .A1(\mem_rdata_q[4] ),
    .S(_20198_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _24095_ (.A0(net58),
    .A1(\mem_rdata_q[3] ),
    .S(_20194_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _24096_ (.A0(net55),
    .A1(\mem_rdata_q[2] ),
    .S(_20194_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _24097_ (.A0(net525),
    .A1(\mem_rdata_q[1] ),
    .S(_20194_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _24098_ (.A0(net33),
    .A1(\mem_rdata_q[0] ),
    .S(_20194_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_1 _24099_ (.A(_19601_),
    .B(_19687_),
    .Y(_20199_));
 sky130_fd_sc_hd__buf_6 _24100_ (.A(_20199_),
    .X(_20200_));
 sky130_fd_sc_hd__clkbuf_4 _24101_ (.A(_20200_),
    .X(_20201_));
 sky130_fd_sc_hd__mux2_1 _24102_ (.A0(_19720_),
    .A1(\cpuregs[18][31] ),
    .S(_20201_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _24103_ (.A0(_19724_),
    .A1(\cpuregs[18][30] ),
    .S(_20201_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _24104_ (.A0(_19725_),
    .A1(\cpuregs[18][29] ),
    .S(_20201_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _24105_ (.A0(_19726_),
    .A1(\cpuregs[18][28] ),
    .S(_20201_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _24106_ (.A0(_19727_),
    .A1(\cpuregs[18][27] ),
    .S(_20201_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _24107_ (.A0(_19728_),
    .A1(\cpuregs[18][26] ),
    .S(_20201_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_4 _24108_ (.A(_20200_),
    .X(_20202_));
 sky130_fd_sc_hd__mux2_1 _24109_ (.A0(_19729_),
    .A1(\cpuregs[18][25] ),
    .S(_20202_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _24110_ (.A0(_19731_),
    .A1(\cpuregs[18][24] ),
    .S(_20202_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _24111_ (.A0(_19732_),
    .A1(\cpuregs[18][23] ),
    .S(_20202_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _24112_ (.A0(_19733_),
    .A1(\cpuregs[18][22] ),
    .S(_20202_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _24113_ (.A0(_19734_),
    .A1(\cpuregs[18][21] ),
    .S(_20202_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _24114_ (.A0(_19735_),
    .A1(\cpuregs[18][20] ),
    .S(_20202_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_4 _24115_ (.A(_20200_),
    .X(_20203_));
 sky130_fd_sc_hd__mux2_1 _24116_ (.A0(_19736_),
    .A1(\cpuregs[18][19] ),
    .S(_20203_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _24117_ (.A0(_19738_),
    .A1(\cpuregs[18][18] ),
    .S(_20203_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _24118_ (.A0(_19739_),
    .A1(\cpuregs[18][17] ),
    .S(_20203_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _24119_ (.A0(_19740_),
    .A1(\cpuregs[18][16] ),
    .S(_20203_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _24120_ (.A0(_19741_),
    .A1(\cpuregs[18][15] ),
    .S(_20203_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _24121_ (.A0(_19742_),
    .A1(\cpuregs[18][14] ),
    .S(_20203_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_4 _24122_ (.A(_20200_),
    .X(_20204_));
 sky130_fd_sc_hd__mux2_1 _24123_ (.A0(_19743_),
    .A1(\cpuregs[18][13] ),
    .S(_20204_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _24124_ (.A0(_19745_),
    .A1(\cpuregs[18][12] ),
    .S(_20204_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _24125_ (.A0(_19746_),
    .A1(\cpuregs[18][11] ),
    .S(_20204_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _24126_ (.A0(_19747_),
    .A1(\cpuregs[18][10] ),
    .S(_20204_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _24127_ (.A0(_19748_),
    .A1(\cpuregs[18][9] ),
    .S(_20204_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _24128_ (.A0(_19749_),
    .A1(\cpuregs[18][8] ),
    .S(_20204_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_4 _24129_ (.A(_20199_),
    .X(_20205_));
 sky130_fd_sc_hd__mux2_1 _24130_ (.A0(_19750_),
    .A1(\cpuregs[18][7] ),
    .S(_20205_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_1 _24131_ (.A0(_19752_),
    .A1(\cpuregs[18][6] ),
    .S(_20205_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _24132_ (.A0(_19753_),
    .A1(\cpuregs[18][5] ),
    .S(_20205_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _24133_ (.A0(_19754_),
    .A1(\cpuregs[18][4] ),
    .S(_20205_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _24134_ (.A0(_19755_),
    .A1(\cpuregs[18][3] ),
    .S(_20205_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _24135_ (.A0(_19756_),
    .A1(\cpuregs[18][2] ),
    .S(_20205_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _24136_ (.A0(_19757_),
    .A1(\cpuregs[18][1] ),
    .S(_20200_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_1 _24137_ (.A0(_19758_),
    .A1(\cpuregs[18][0] ),
    .S(_20200_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_1 _24138_ (.A(_19601_),
    .B(_19644_),
    .Y(_20206_));
 sky130_fd_sc_hd__buf_6 _24139_ (.A(_20206_),
    .X(_20207_));
 sky130_fd_sc_hd__clkbuf_4 _24140_ (.A(_20207_),
    .X(_20208_));
 sky130_fd_sc_hd__mux2_1 _24141_ (.A0(_19767_),
    .A1(\cpuregs[10][31] ),
    .S(_20208_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _24142_ (.A0(_19771_),
    .A1(\cpuregs[10][30] ),
    .S(_20208_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _24143_ (.A0(_19772_),
    .A1(\cpuregs[10][29] ),
    .S(_20208_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _24144_ (.A0(_19773_),
    .A1(\cpuregs[10][28] ),
    .S(_20208_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _24145_ (.A0(_19774_),
    .A1(\cpuregs[10][27] ),
    .S(_20208_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _24146_ (.A0(_19775_),
    .A1(\cpuregs[10][26] ),
    .S(_20208_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_4 _24147_ (.A(_20207_),
    .X(_20209_));
 sky130_fd_sc_hd__mux2_1 _24148_ (.A0(_19776_),
    .A1(\cpuregs[10][25] ),
    .S(_20209_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _24149_ (.A0(_19778_),
    .A1(\cpuregs[10][24] ),
    .S(_20209_),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_1 _24150_ (.A0(_19779_),
    .A1(\cpuregs[10][23] ),
    .S(_20209_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _24151_ (.A0(_19780_),
    .A1(\cpuregs[10][22] ),
    .S(_20209_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _24152_ (.A0(_19781_),
    .A1(\cpuregs[10][21] ),
    .S(_20209_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _24153_ (.A0(_19782_),
    .A1(\cpuregs[10][20] ),
    .S(_20209_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_4 _24154_ (.A(_20207_),
    .X(_20210_));
 sky130_fd_sc_hd__mux2_1 _24155_ (.A0(_19783_),
    .A1(\cpuregs[10][19] ),
    .S(_20210_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _24156_ (.A0(_19785_),
    .A1(\cpuregs[10][18] ),
    .S(_20210_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _24157_ (.A0(_19786_),
    .A1(\cpuregs[10][17] ),
    .S(_20210_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _24158_ (.A0(_19787_),
    .A1(\cpuregs[10][16] ),
    .S(_20210_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _24159_ (.A0(_19788_),
    .A1(\cpuregs[10][15] ),
    .S(_20210_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _24160_ (.A0(_19789_),
    .A1(\cpuregs[10][14] ),
    .S(_20210_),
    .X(_02881_));
 sky130_fd_sc_hd__buf_4 _24161_ (.A(_20207_),
    .X(_20211_));
 sky130_fd_sc_hd__mux2_1 _24162_ (.A0(_19790_),
    .A1(\cpuregs[10][13] ),
    .S(_20211_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _24163_ (.A0(_19792_),
    .A1(\cpuregs[10][12] ),
    .S(_20211_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _24164_ (.A0(_19793_),
    .A1(\cpuregs[10][11] ),
    .S(_20211_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _24165_ (.A0(_19794_),
    .A1(\cpuregs[10][10] ),
    .S(_20211_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _24166_ (.A0(_19795_),
    .A1(\cpuregs[10][9] ),
    .S(_20211_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _24167_ (.A0(_19796_),
    .A1(\cpuregs[10][8] ),
    .S(_20211_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_4 _24168_ (.A(_20206_),
    .X(_20212_));
 sky130_fd_sc_hd__mux2_1 _24169_ (.A0(_19797_),
    .A1(\cpuregs[10][7] ),
    .S(_20212_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _24170_ (.A0(_19799_),
    .A1(\cpuregs[10][6] ),
    .S(_20212_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _24171_ (.A0(_19800_),
    .A1(\cpuregs[10][5] ),
    .S(_20212_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _24172_ (.A0(_19801_),
    .A1(\cpuregs[10][4] ),
    .S(_20212_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _24173_ (.A0(_19802_),
    .A1(\cpuregs[10][3] ),
    .S(_20212_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _24174_ (.A0(_19803_),
    .A1(\cpuregs[10][2] ),
    .S(_20212_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _24175_ (.A0(_19804_),
    .A1(\cpuregs[10][1] ),
    .S(_20207_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _24176_ (.A0(_19805_),
    .A1(\cpuregs[10][0] ),
    .S(_20207_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _24177_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _24178_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _24179_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _24180_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _24181_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _24182_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _24183_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _24184_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _24185_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _24186_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _24187_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _24188_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _24189_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _24190_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _24191_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _24192_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _24193_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _24194_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _24195_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _24196_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _24197_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _24198_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _24199_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _24200_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _24201_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _24202_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _24203_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _24204_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _24205_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _24206_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _24207_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _24208_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_1 _24209_ (.A(_19601_),
    .B(_19712_),
    .Y(_20213_));
 sky130_fd_sc_hd__buf_6 _24210_ (.A(_20213_),
    .X(_20214_));
 sky130_fd_sc_hd__clkbuf_4 _24211_ (.A(_20214_),
    .X(_20215_));
 sky130_fd_sc_hd__mux2_1 _24212_ (.A0(_19767_),
    .A1(\cpuregs[14][31] ),
    .S(_20215_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _24213_ (.A0(_19771_),
    .A1(\cpuregs[14][30] ),
    .S(_20215_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _24214_ (.A0(_19772_),
    .A1(\cpuregs[14][29] ),
    .S(_20215_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _24215_ (.A0(_19773_),
    .A1(\cpuregs[14][28] ),
    .S(_20215_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _24216_ (.A0(_19774_),
    .A1(\cpuregs[14][27] ),
    .S(_20215_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _24217_ (.A0(_19775_),
    .A1(\cpuregs[14][26] ),
    .S(_20215_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_4 _24218_ (.A(_20214_),
    .X(_20216_));
 sky130_fd_sc_hd__mux2_1 _24219_ (.A0(_19776_),
    .A1(\cpuregs[14][25] ),
    .S(_20216_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _24220_ (.A0(_19778_),
    .A1(\cpuregs[14][24] ),
    .S(_20216_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _24221_ (.A0(_19779_),
    .A1(\cpuregs[14][23] ),
    .S(_20216_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _24222_ (.A0(_19780_),
    .A1(\cpuregs[14][22] ),
    .S(_20216_),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_1 _24223_ (.A0(_19781_),
    .A1(\cpuregs[14][21] ),
    .S(_20216_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _24224_ (.A0(_19782_),
    .A1(\cpuregs[14][20] ),
    .S(_20216_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_4 _24225_ (.A(_20214_),
    .X(_20217_));
 sky130_fd_sc_hd__mux2_1 _24226_ (.A0(_19783_),
    .A1(\cpuregs[14][19] ),
    .S(_20217_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _24227_ (.A0(_19785_),
    .A1(\cpuregs[14][18] ),
    .S(_20217_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _24228_ (.A0(_19786_),
    .A1(\cpuregs[14][17] ),
    .S(_20217_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _24229_ (.A0(_19787_),
    .A1(\cpuregs[14][16] ),
    .S(_20217_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _24230_ (.A0(_19788_),
    .A1(\cpuregs[14][15] ),
    .S(_20217_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _24231_ (.A0(_19789_),
    .A1(\cpuregs[14][14] ),
    .S(_20217_),
    .X(_02817_));
 sky130_fd_sc_hd__buf_4 _24232_ (.A(_20214_),
    .X(_20218_));
 sky130_fd_sc_hd__mux2_1 _24233_ (.A0(_19790_),
    .A1(\cpuregs[14][13] ),
    .S(_20218_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _24234_ (.A0(_19792_),
    .A1(\cpuregs[14][12] ),
    .S(_20218_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _24235_ (.A0(_19793_),
    .A1(\cpuregs[14][11] ),
    .S(_20218_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _24236_ (.A0(_19794_),
    .A1(\cpuregs[14][10] ),
    .S(_20218_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _24237_ (.A0(_19795_),
    .A1(\cpuregs[14][9] ),
    .S(_20218_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _24238_ (.A0(_19796_),
    .A1(\cpuregs[14][8] ),
    .S(_20218_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_4 _24239_ (.A(_20213_),
    .X(_20219_));
 sky130_fd_sc_hd__mux2_1 _24240_ (.A0(_19797_),
    .A1(\cpuregs[14][7] ),
    .S(_20219_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _24241_ (.A0(_19799_),
    .A1(\cpuregs[14][6] ),
    .S(_20219_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _24242_ (.A0(_19800_),
    .A1(\cpuregs[14][5] ),
    .S(_20219_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _24243_ (.A0(_19801_),
    .A1(\cpuregs[14][4] ),
    .S(_20219_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _24244_ (.A0(_19802_),
    .A1(\cpuregs[14][3] ),
    .S(_20219_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _24245_ (.A0(_19803_),
    .A1(\cpuregs[14][2] ),
    .S(_20219_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _24246_ (.A0(_19804_),
    .A1(\cpuregs[14][1] ),
    .S(_20214_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _24247_ (.A0(_19805_),
    .A1(\cpuregs[14][0] ),
    .S(_20214_),
    .X(_02803_));
 sky130_fd_sc_hd__or3_1 _24248_ (.A(_19592_),
    .B(_19643_),
    .C(_19599_),
    .X(_20220_));
 sky130_fd_sc_hd__buf_6 _24249_ (.A(_20220_),
    .X(_20221_));
 sky130_fd_sc_hd__buf_4 _24250_ (.A(_20221_),
    .X(_20222_));
 sky130_fd_sc_hd__mux2_1 _24251_ (.A0(_19767_),
    .A1(\cpuregs[8][31] ),
    .S(_20222_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _24252_ (.A0(_19771_),
    .A1(\cpuregs[8][30] ),
    .S(_20222_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _24253_ (.A0(_19772_),
    .A1(\cpuregs[8][29] ),
    .S(_20222_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _24254_ (.A0(_19773_),
    .A1(\cpuregs[8][28] ),
    .S(_20222_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _24255_ (.A0(_19774_),
    .A1(\cpuregs[8][27] ),
    .S(_20222_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _24256_ (.A0(_19775_),
    .A1(\cpuregs[8][26] ),
    .S(_20222_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_4 _24257_ (.A(_20221_),
    .X(_20223_));
 sky130_fd_sc_hd__mux2_1 _24258_ (.A0(_19776_),
    .A1(\cpuregs[8][25] ),
    .S(_20223_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _24259_ (.A0(_19778_),
    .A1(\cpuregs[8][24] ),
    .S(_20223_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _24260_ (.A0(_19779_),
    .A1(\cpuregs[8][23] ),
    .S(_20223_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _24261_ (.A0(_19780_),
    .A1(\cpuregs[8][22] ),
    .S(_20223_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _24262_ (.A0(_19781_),
    .A1(\cpuregs[8][21] ),
    .S(_20223_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _24263_ (.A0(_19782_),
    .A1(\cpuregs[8][20] ),
    .S(_20223_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_4 _24264_ (.A(_20221_),
    .X(_20224_));
 sky130_fd_sc_hd__mux2_1 _24265_ (.A0(_19783_),
    .A1(\cpuregs[8][19] ),
    .S(_20224_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _24266_ (.A0(_19785_),
    .A1(\cpuregs[8][18] ),
    .S(_20224_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _24267_ (.A0(_19786_),
    .A1(\cpuregs[8][17] ),
    .S(_20224_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_1 _24268_ (.A0(_19787_),
    .A1(\cpuregs[8][16] ),
    .S(_20224_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _24269_ (.A0(_19788_),
    .A1(\cpuregs[8][15] ),
    .S(_20224_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _24270_ (.A0(_19789_),
    .A1(\cpuregs[8][14] ),
    .S(_20224_),
    .X(_02785_));
 sky130_fd_sc_hd__buf_4 _24271_ (.A(_20221_),
    .X(_20225_));
 sky130_fd_sc_hd__mux2_1 _24272_ (.A0(_19790_),
    .A1(\cpuregs[8][13] ),
    .S(_20225_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _24273_ (.A0(_19792_),
    .A1(\cpuregs[8][12] ),
    .S(_20225_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _24274_ (.A0(_19793_),
    .A1(\cpuregs[8][11] ),
    .S(_20225_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _24275_ (.A0(_19794_),
    .A1(\cpuregs[8][10] ),
    .S(_20225_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _24276_ (.A0(_19795_),
    .A1(\cpuregs[8][9] ),
    .S(_20225_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _24277_ (.A0(_19796_),
    .A1(\cpuregs[8][8] ),
    .S(_20225_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_4 _24278_ (.A(_20220_),
    .X(_20226_));
 sky130_fd_sc_hd__mux2_1 _24279_ (.A0(_19797_),
    .A1(\cpuregs[8][7] ),
    .S(_20226_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _24280_ (.A0(_19799_),
    .A1(\cpuregs[8][6] ),
    .S(_20226_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _24281_ (.A0(_19800_),
    .A1(\cpuregs[8][5] ),
    .S(_20226_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _24282_ (.A0(_19801_),
    .A1(\cpuregs[8][4] ),
    .S(_20226_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _24283_ (.A0(_19802_),
    .A1(\cpuregs[8][3] ),
    .S(_20226_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _24284_ (.A0(_19803_),
    .A1(\cpuregs[8][2] ),
    .S(_20226_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _24285_ (.A0(_19804_),
    .A1(\cpuregs[8][1] ),
    .S(_20221_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _24286_ (.A0(_19805_),
    .A1(\cpuregs[8][0] ),
    .S(_20221_),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_8 _24287_ (.A(latched_branch),
    .B(_18748_),
    .Y(_00292_));
 sky130_fd_sc_hd__nor2_1 _24288_ (.A(latched_store),
    .B(_18555_),
    .Y(_20227_));
 sky130_fd_sc_hd__o311a_1 _24289_ (.A1(_18967_),
    .A2(net472),
    .A3(_20227_),
    .B1(_18543_),
    .C1(\reg_next_pc[0] ),
    .X(_02770_));
 sky130_fd_sc_hd__and2_1 _24290_ (.A(_19403_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_1 _24291_ (.A(_19403_),
    .B(_21143_),
    .X(_02768_));
 sky130_fd_sc_hd__and2_1 _24292_ (.A(_19403_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__clkbuf_2 _24293_ (.A(_19399_),
    .X(_20228_));
 sky130_fd_sc_hd__and2_1 _24294_ (.A(_20228_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _24295_ (.A(_20228_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_1 _24296_ (.A(_20228_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_1 _24297_ (.A(_20228_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__and2_1 _24298_ (.A(_20228_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__and2_1 _24299_ (.A(_20228_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_2 _24300_ (.A(_19399_),
    .X(_20229_));
 sky130_fd_sc_hd__and2_1 _24301_ (.A(_20229_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__and2_1 _24302_ (.A(_20229_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_1 _24303_ (.A(_20229_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_1 _24304_ (.A(_20229_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_1 _24305_ (.A(_20229_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_1 _24306_ (.A(_20229_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__buf_1 _24307_ (.A(_18548_),
    .X(_20230_));
 sky130_fd_sc_hd__and2_1 _24308_ (.A(_20230_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_1 _24309_ (.A(_20230_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_1 _24310_ (.A(_20230_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_1 _24311_ (.A(_20230_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__and2_1 _24312_ (.A(_20230_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_1 _24313_ (.A(_20230_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_2 _24314_ (.A(_18548_),
    .X(_20231_));
 sky130_fd_sc_hd__and2_1 _24315_ (.A(_20231_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_1 _24316_ (.A(_20231_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_1 _24317_ (.A(_20231_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_1 _24318_ (.A(_20231_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_1 _24319_ (.A(_20231_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_1 _24320_ (.A(_20231_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_1 _24321_ (.A(_18703_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_1 _24322_ (.A(_18703_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_1 _24323_ (.A(_18703_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_1 _24324_ (.A(_18703_),
    .B(_00030_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_1 _24325_ (.A(_19972_),
    .B(\mem_rdata_q[21] ),
    .Y(_20232_));
 sky130_fd_sc_hd__clkbuf_2 _24326_ (.A(instr_jal),
    .X(_20233_));
 sky130_fd_sc_hd__clkbuf_2 _24327_ (.A(_20233_),
    .X(_20234_));
 sky130_fd_sc_hd__nand2_1 _24328_ (.A(\decoded_imm_uj[1] ),
    .B(_20234_),
    .Y(_20235_));
 sky130_fd_sc_hd__nor2_1 _24329_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(is_sb_sh_sw),
    .Y(_20236_));
 sky130_fd_sc_hd__inv_2 _24330_ (.A(_20236_),
    .Y(_20237_));
 sky130_fd_sc_hd__nand2_1 _24331_ (.A(_20237_),
    .B(\mem_rdata_q[8] ),
    .Y(_20238_));
 sky130_fd_sc_hd__a31o_1 _24332_ (.A1(_20232_),
    .A2(_20235_),
    .A3(_20238_),
    .B1(_18908_),
    .X(_20239_));
 sky130_fd_sc_hd__a21bo_1 _24333_ (.A1(\decoded_imm[1] ),
    .A2(_20007_),
    .B1_N(_20239_),
    .X(_02738_));
 sky130_vsdinv _24334_ (.A(\decoded_imm[2] ),
    .Y(_20240_));
 sky130_fd_sc_hd__nand2_1 _24335_ (.A(_19972_),
    .B(\mem_rdata_q[22] ),
    .Y(_20241_));
 sky130_fd_sc_hd__nand2_1 _24336_ (.A(\decoded_imm_uj[2] ),
    .B(_18782_),
    .Y(_20242_));
 sky130_fd_sc_hd__nand2_1 _24337_ (.A(_20237_),
    .B(\mem_rdata_q[9] ),
    .Y(_20243_));
 sky130_fd_sc_hd__a31o_1 _24338_ (.A1(_20241_),
    .A2(_20242_),
    .A3(_20243_),
    .B1(_18871_),
    .X(_20244_));
 sky130_fd_sc_hd__o21ai_1 _24339_ (.A1(_20240_),
    .A2(_19955_),
    .B1(_20244_),
    .Y(_02737_));
 sky130_fd_sc_hd__nand2_1 _24340_ (.A(_19972_),
    .B(\mem_rdata_q[23] ),
    .Y(_20245_));
 sky130_fd_sc_hd__clkbuf_2 _24341_ (.A(_20233_),
    .X(_20246_));
 sky130_fd_sc_hd__nand2_1 _24342_ (.A(\decoded_imm_uj[3] ),
    .B(_20246_),
    .Y(_20247_));
 sky130_fd_sc_hd__nand2_1 _24343_ (.A(_20237_),
    .B(\mem_rdata_q[10] ),
    .Y(_20248_));
 sky130_fd_sc_hd__a31o_1 _24344_ (.A1(_20245_),
    .A2(_20247_),
    .A3(_20248_),
    .B1(_18908_),
    .X(_20249_));
 sky130_fd_sc_hd__a21bo_1 _24345_ (.A1(\decoded_imm[3] ),
    .A2(_20007_),
    .B1_N(_20249_),
    .X(_02736_));
 sky130_vsdinv _24346_ (.A(\decoded_imm[4] ),
    .Y(_20250_));
 sky130_fd_sc_hd__nand2_1 _24347_ (.A(_19972_),
    .B(\mem_rdata_q[24] ),
    .Y(_20251_));
 sky130_fd_sc_hd__nand2_1 _24348_ (.A(\decoded_imm_uj[4] ),
    .B(_18782_),
    .Y(_20252_));
 sky130_fd_sc_hd__nand2_1 _24349_ (.A(_20237_),
    .B(\mem_rdata_q[11] ),
    .Y(_20253_));
 sky130_fd_sc_hd__a31o_1 _24350_ (.A1(_20251_),
    .A2(_20252_),
    .A3(_20253_),
    .B1(_18871_),
    .X(_20254_));
 sky130_fd_sc_hd__o21ai_1 _24351_ (.A1(_20250_),
    .A2(_19955_),
    .B1(_20254_),
    .Y(_02735_));
 sky130_fd_sc_hd__nor2_2 _24352_ (.A(_20237_),
    .B(_19971_),
    .Y(_20255_));
 sky130_vsdinv _24353_ (.A(_20255_),
    .Y(_20256_));
 sky130_fd_sc_hd__a22o_1 _24354_ (.A1(\decoded_imm_uj[5] ),
    .A2(_18782_),
    .B1(_20256_),
    .B2(_18898_),
    .X(_20257_));
 sky130_fd_sc_hd__mux2_1 _24355_ (.A0(_20257_),
    .A1(\decoded_imm[5] ),
    .S(_18905_),
    .X(_02734_));
 sky130_fd_sc_hd__a22o_1 _24356_ (.A1(\decoded_imm_uj[6] ),
    .A2(_18782_),
    .B1(_20256_),
    .B2(\mem_rdata_q[26] ),
    .X(_20258_));
 sky130_fd_sc_hd__mux2_1 _24357_ (.A0(_20258_),
    .A1(\decoded_imm[6] ),
    .S(_18905_),
    .X(_02733_));
 sky130_fd_sc_hd__a22o_1 _24358_ (.A1(\decoded_imm_uj[7] ),
    .A2(_20234_),
    .B1(_20256_),
    .B2(\mem_rdata_q[27] ),
    .X(_20259_));
 sky130_fd_sc_hd__buf_2 _24359_ (.A(_18904_),
    .X(_20260_));
 sky130_fd_sc_hd__mux2_1 _24360_ (.A0(_20259_),
    .A1(\decoded_imm[7] ),
    .S(_20260_),
    .X(_02732_));
 sky130_fd_sc_hd__a22o_1 _24361_ (.A1(\decoded_imm_uj[8] ),
    .A2(_20234_),
    .B1(_20256_),
    .B2(\mem_rdata_q[28] ),
    .X(_20261_));
 sky130_fd_sc_hd__mux2_1 _24362_ (.A0(_20261_),
    .A1(\decoded_imm[8] ),
    .S(_20260_),
    .X(_02731_));
 sky130_fd_sc_hd__a22o_1 _24363_ (.A1(\decoded_imm_uj[9] ),
    .A2(_20234_),
    .B1(_20256_),
    .B2(\mem_rdata_q[29] ),
    .X(_20262_));
 sky130_fd_sc_hd__mux2_1 _24364_ (.A0(_20262_),
    .A1(\decoded_imm[9] ),
    .S(_20260_),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_1 _24365_ (.A1(\decoded_imm_uj[10] ),
    .A2(_20234_),
    .B1(_20256_),
    .B2(\mem_rdata_q[30] ),
    .X(_20263_));
 sky130_fd_sc_hd__mux2_1 _24366_ (.A0(_20263_),
    .A1(\decoded_imm[10] ),
    .S(_20260_),
    .X(_02729_));
 sky130_fd_sc_hd__o21a_1 _24367_ (.A1(_19951_),
    .A2(_19971_),
    .B1(_20024_),
    .X(_20264_));
 sky130_fd_sc_hd__a221o_1 _24368_ (.A1(_18699_),
    .A2(\mem_rdata_q[7] ),
    .B1(\decoded_imm_uj[11] ),
    .B2(_20233_),
    .C1(_20264_),
    .X(_20265_));
 sky130_fd_sc_hd__mux2_1 _24369_ (.A0(_20265_),
    .A1(\decoded_imm[11] ),
    .S(_20260_),
    .X(_02728_));
 sky130_vsdinv _24370_ (.A(_18737_),
    .Y(_20266_));
 sky130_fd_sc_hd__clkbuf_2 _24371_ (.A(_20266_),
    .X(_20267_));
 sky130_fd_sc_hd__nor2_2 _24372_ (.A(_18876_),
    .B(_20255_),
    .Y(_20268_));
 sky130_fd_sc_hd__clkbuf_2 _24373_ (.A(_20268_),
    .X(_20269_));
 sky130_fd_sc_hd__a221o_1 _24374_ (.A1(\decoded_imm_uj[12] ),
    .A2(_20246_),
    .B1(_18889_),
    .B2(_20267_),
    .C1(_20269_),
    .X(_20270_));
 sky130_fd_sc_hd__mux2_1 _24375_ (.A0(_20270_),
    .A1(\decoded_imm[12] ),
    .S(_20260_),
    .X(_02727_));
 sky130_fd_sc_hd__a221o_1 _24376_ (.A1(\decoded_imm_uj[13] ),
    .A2(_20246_),
    .B1(\mem_rdata_q[13] ),
    .B2(_20267_),
    .C1(_20269_),
    .X(_20271_));
 sky130_fd_sc_hd__buf_2 _24377_ (.A(_18870_),
    .X(_20272_));
 sky130_fd_sc_hd__mux2_1 _24378_ (.A0(_20271_),
    .A1(\decoded_imm[13] ),
    .S(_20272_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_2 _24379_ (.A(_20266_),
    .X(_20273_));
 sky130_fd_sc_hd__a221o_1 _24380_ (.A1(\decoded_imm_uj[14] ),
    .A2(_20246_),
    .B1(_18893_),
    .B2(_20273_),
    .C1(_20269_),
    .X(_20274_));
 sky130_fd_sc_hd__mux2_1 _24381_ (.A0(_20274_),
    .A1(\decoded_imm[14] ),
    .S(_20272_),
    .X(_02725_));
 sky130_fd_sc_hd__a221o_1 _24382_ (.A1(\decoded_imm_uj[15] ),
    .A2(_20246_),
    .B1(\mem_rdata_q[15] ),
    .B2(_20273_),
    .C1(_20269_),
    .X(_20275_));
 sky130_fd_sc_hd__mux2_1 _24383_ (.A0(_20275_),
    .A1(\decoded_imm[15] ),
    .S(_20272_),
    .X(_02724_));
 sky130_fd_sc_hd__a221o_1 _24384_ (.A1(\decoded_imm_uj[16] ),
    .A2(_20246_),
    .B1(\mem_rdata_q[16] ),
    .B2(_20273_),
    .C1(_20269_),
    .X(_20276_));
 sky130_fd_sc_hd__mux2_1 _24385_ (.A0(_20276_),
    .A1(\decoded_imm[16] ),
    .S(_20272_),
    .X(_02723_));
 sky130_fd_sc_hd__a221o_1 _24386_ (.A1(\decoded_imm_uj[17] ),
    .A2(_20233_),
    .B1(\mem_rdata_q[17] ),
    .B2(_20273_),
    .C1(_20269_),
    .X(_20277_));
 sky130_fd_sc_hd__mux2_1 _24387_ (.A0(_20277_),
    .A1(\decoded_imm[17] ),
    .S(_20272_),
    .X(_02722_));
 sky130_fd_sc_hd__a221o_1 _24388_ (.A1(\decoded_imm_uj[18] ),
    .A2(_20233_),
    .B1(\mem_rdata_q[18] ),
    .B2(_20273_),
    .C1(_20268_),
    .X(_20278_));
 sky130_fd_sc_hd__mux2_1 _24389_ (.A0(_20278_),
    .A1(\decoded_imm[18] ),
    .S(_20272_),
    .X(_02721_));
 sky130_fd_sc_hd__a221o_1 _24390_ (.A1(\decoded_imm_uj[19] ),
    .A2(_20233_),
    .B1(\mem_rdata_q[19] ),
    .B2(_20273_),
    .C1(_20268_),
    .X(_20279_));
 sky130_fd_sc_hd__mux2_1 _24391_ (.A0(_20279_),
    .A1(\decoded_imm[19] ),
    .S(_18871_),
    .X(_02720_));
 sky130_fd_sc_hd__a22o_2 _24392_ (.A1(_19961_),
    .A2(instr_jal),
    .B1(_20237_),
    .B2(_20024_),
    .X(_20280_));
 sky130_fd_sc_hd__clkbuf_2 _24393_ (.A(_20280_),
    .X(_20281_));
 sky130_fd_sc_hd__and2_2 _24394_ (.A(_19972_),
    .B(_20024_),
    .X(_20282_));
 sky130_fd_sc_hd__a21o_1 _24395_ (.A1(\mem_rdata_q[20] ),
    .A2(_20267_),
    .B1(_18930_),
    .X(_20283_));
 sky130_fd_sc_hd__o32a_1 _24396_ (.A1(_20281_),
    .A2(_20282_),
    .A3(_20283_),
    .B1(\decoded_imm[20] ),
    .B2(_19955_),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_2 _24397_ (.A(_18737_),
    .X(_20284_));
 sky130_fd_sc_hd__o21ai_1 _24398_ (.A1(_20002_),
    .A2(_20284_),
    .B1(_20030_),
    .Y(_20285_));
 sky130_fd_sc_hd__clkbuf_2 _24399_ (.A(_20282_),
    .X(_20286_));
 sky130_fd_sc_hd__o32a_1 _24400_ (.A1(_20285_),
    .A2(_20281_),
    .A3(_20286_),
    .B1(\decoded_imm[21] ),
    .B2(_19955_),
    .X(_02718_));
 sky130_fd_sc_hd__a21o_1 _24401_ (.A1(\mem_rdata_q[22] ),
    .A2(_20267_),
    .B1(_18904_),
    .X(_20287_));
 sky130_fd_sc_hd__clkbuf_2 _24402_ (.A(_18922_),
    .X(_20288_));
 sky130_fd_sc_hd__o32a_1 _24403_ (.A1(_20281_),
    .A2(_20282_),
    .A3(_20287_),
    .B1(\decoded_imm[22] ),
    .B2(_20288_),
    .X(_02717_));
 sky130_fd_sc_hd__a21o_1 _24404_ (.A1(\mem_rdata_q[23] ),
    .A2(_20267_),
    .B1(_18904_),
    .X(_20289_));
 sky130_fd_sc_hd__o32a_1 _24405_ (.A1(_20281_),
    .A2(_20282_),
    .A3(_20289_),
    .B1(\decoded_imm[23] ),
    .B2(_20288_),
    .X(_02716_));
 sky130_fd_sc_hd__o21ai_1 _24406_ (.A1(_19997_),
    .A2(_20284_),
    .B1(_20030_),
    .Y(_20290_));
 sky130_fd_sc_hd__o32a_1 _24407_ (.A1(_20290_),
    .A2(_20281_),
    .A3(_20286_),
    .B1(\decoded_imm[24] ),
    .B2(_20288_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ai_1 _24408_ (.A1(_18884_),
    .A2(_20284_),
    .B1(_18918_),
    .Y(_20291_));
 sky130_fd_sc_hd__o32a_1 _24409_ (.A1(_20291_),
    .A2(_20280_),
    .A3(_20286_),
    .B1(\decoded_imm[25] ),
    .B2(_20288_),
    .X(_02714_));
 sky130_fd_sc_hd__a21o_1 _24410_ (.A1(\mem_rdata_q[26] ),
    .A2(_20267_),
    .B1(_18904_),
    .X(_20292_));
 sky130_fd_sc_hd__o32a_1 _24411_ (.A1(_20281_),
    .A2(_20282_),
    .A3(_20292_),
    .B1(\decoded_imm[26] ),
    .B2(_20288_),
    .X(_02713_));
 sky130_fd_sc_hd__o21ai_1 _24412_ (.A1(_18880_),
    .A2(_20284_),
    .B1(_18918_),
    .Y(_20293_));
 sky130_fd_sc_hd__o32a_1 _24413_ (.A1(_20293_),
    .A2(_20280_),
    .A3(_20286_),
    .B1(\decoded_imm[27] ),
    .B2(_20288_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_1 _24414_ (.A1(_19983_),
    .A2(_20284_),
    .B1(_18918_),
    .Y(_20294_));
 sky130_fd_sc_hd__o32a_1 _24415_ (.A1(_20294_),
    .A2(_20280_),
    .A3(_20286_),
    .B1(\decoded_imm[28] ),
    .B2(_20025_),
    .X(_02711_));
 sky130_fd_sc_hd__o21ai_1 _24416_ (.A1(_18878_),
    .A2(_20284_),
    .B1(_18918_),
    .Y(_20295_));
 sky130_fd_sc_hd__o32a_1 _24417_ (.A1(_20295_),
    .A2(_20280_),
    .A3(_20286_),
    .B1(\decoded_imm[29] ),
    .B2(_20025_),
    .X(_02710_));
 sky130_fd_sc_hd__o21ai_1 _24418_ (.A1(_18877_),
    .A2(_18737_),
    .B1(_18918_),
    .Y(_20296_));
 sky130_fd_sc_hd__o32a_1 _24419_ (.A1(_20296_),
    .A2(_20280_),
    .A3(_20282_),
    .B1(\decoded_imm[30] ),
    .B2(_20025_),
    .X(_02709_));
 sky130_fd_sc_hd__nand2_1 _24420_ (.A(_20255_),
    .B(_18737_),
    .Y(_20297_));
 sky130_fd_sc_hd__a22o_1 _24421_ (.A1(_19962_),
    .A2(_20234_),
    .B1(_20297_),
    .B2(_20024_),
    .X(_20298_));
 sky130_fd_sc_hd__mux2_1 _24422_ (.A0(_20298_),
    .A1(\decoded_imm[31] ),
    .S(_18871_),
    .X(_02708_));
 sky130_fd_sc_hd__and4_4 _24423_ (.A(_19710_),
    .B(_18540_),
    .C(_18706_),
    .D(_18553_),
    .X(_20299_));
 sky130_fd_sc_hd__clkbuf_2 _24424_ (.A(_20299_),
    .X(_20300_));
 sky130_fd_sc_hd__nor2_1 _24425_ (.A(_19591_),
    .B(_20300_),
    .Y(_20301_));
 sky130_fd_sc_hd__a31o_1 _24426_ (.A1(_21103_),
    .A2(_18719_),
    .A3(_20300_),
    .B1(_20301_),
    .X(_02707_));
 sky130_fd_sc_hd__nor2_8 _24427_ (.A(_02542_),
    .B(net414),
    .Y(_20302_));
 sky130_fd_sc_hd__nor2_1 _24428_ (.A(_19590_),
    .B(_20300_),
    .Y(_20303_));
 sky130_fd_sc_hd__a31o_1 _24429_ (.A1(_20302_),
    .A2(\decoded_rd[1] ),
    .A3(_20300_),
    .B1(_20303_),
    .X(_02706_));
 sky130_fd_sc_hd__nor2_1 _24430_ (.A(_19686_),
    .B(_20299_),
    .Y(_20304_));
 sky130_fd_sc_hd__a31o_1 _24431_ (.A1(_20302_),
    .A2(\decoded_rd[2] ),
    .A3(_20300_),
    .B1(_20304_),
    .X(_02705_));
 sky130_fd_sc_hd__nor2_1 _24432_ (.A(_19594_),
    .B(_20299_),
    .Y(_20305_));
 sky130_fd_sc_hd__a31o_1 _24433_ (.A1(_20302_),
    .A2(\decoded_rd[3] ),
    .A3(_20300_),
    .B1(_20305_),
    .X(_02704_));
 sky130_fd_sc_hd__nor2_4 _24434_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .Y(_01304_));
 sky130_vsdinv _24435_ (.A(is_lui_auipc_jal),
    .Y(_20306_));
 sky130_fd_sc_hd__a21o_1 _24436_ (.A1(_01304_),
    .A2(_20306_),
    .B1(_19316_),
    .X(_20307_));
 sky130_fd_sc_hd__o31a_1 _24437_ (.A1(_19951_),
    .A2(_18743_),
    .A3(_00310_),
    .B1(_20307_),
    .X(_20308_));
 sky130_fd_sc_hd__nor2b_1 _24438_ (.A(_20308_),
    .B_N(_19654_),
    .Y(_02703_));
 sky130_vsdinv _24439_ (.A(net226),
    .Y(_20309_));
 sky130_fd_sc_hd__clkbuf_2 _24440_ (.A(_20309_),
    .X(_20310_));
 sky130_fd_sc_hd__clkbuf_2 _24441_ (.A(_20310_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_1 _24442_ (.A(_02327_),
    .B(_02558_),
    .X(_02702_));
 sky130_fd_sc_hd__and2_1 _24443_ (.A(_02327_),
    .B(_02557_),
    .X(_02701_));
 sky130_fd_sc_hd__and2_1 _24444_ (.A(_02327_),
    .B(_02556_),
    .X(_02700_));
 sky130_fd_sc_hd__and2_1 _24445_ (.A(_02327_),
    .B(_02555_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_1 _24446_ (.A(_20310_),
    .B(_02554_),
    .X(_02698_));
 sky130_fd_sc_hd__and2_1 _24447_ (.A(_20310_),
    .B(_02553_),
    .X(_02697_));
 sky130_fd_sc_hd__and2_1 _24448_ (.A(_20310_),
    .B(_02552_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_1 _24449_ (.A(_20310_),
    .B(_02551_),
    .X(_02695_));
 sky130_fd_sc_hd__clkbuf_4 _24450_ (.A(_19674_),
    .X(_20311_));
 sky130_vsdinv _24451_ (.A(_00122_),
    .Y(_20312_));
 sky130_fd_sc_hd__nor2_1 _24452_ (.A(_20311_),
    .B(_20312_),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_2 _24453_ (.A(_19673_),
    .B(_19674_),
    .Y(_20313_));
 sky130_vsdinv _24454_ (.A(_20313_),
    .Y(_20314_));
 sky130_fd_sc_hd__nor2_1 _24455_ (.A(_20312_),
    .B(_20314_),
    .Y(_02694_));
 sky130_vsdinv _24456_ (.A(_00116_),
    .Y(_20315_));
 sky130_fd_sc_hd__nor2_1 _24457_ (.A(_20311_),
    .B(_20315_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor2_1 _24458_ (.A(_20315_),
    .B(_20314_),
    .Y(_02693_));
 sky130_vsdinv _24459_ (.A(_00110_),
    .Y(_20316_));
 sky130_fd_sc_hd__nor2_1 _24460_ (.A(_20311_),
    .B(_20316_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor2_1 _24461_ (.A(_20316_),
    .B(_20314_),
    .Y(_02692_));
 sky130_vsdinv _24462_ (.A(_00104_),
    .Y(_20317_));
 sky130_fd_sc_hd__nor2_1 _24463_ (.A(_20311_),
    .B(_20317_),
    .Y(_02547_));
 sky130_fd_sc_hd__nor2_1 _24464_ (.A(_20317_),
    .B(_20314_),
    .Y(_02691_));
 sky130_fd_sc_hd__nor2_4 _24465_ (.A(net225),
    .B(net222),
    .Y(_20318_));
 sky130_fd_sc_hd__and2_1 _24466_ (.A(_20318_),
    .B(_00094_),
    .X(_02546_));
 sky130_vsdinv _24467_ (.A(net222),
    .Y(_20319_));
 sky130_fd_sc_hd__clkbuf_2 _24468_ (.A(_20319_),
    .X(_02321_));
 sky130_fd_sc_hd__and3_1 _24469_ (.A(_20313_),
    .B(_02321_),
    .C(_00094_),
    .X(_02690_));
 sky130_fd_sc_hd__and2_1 _24470_ (.A(_20318_),
    .B(_00084_),
    .X(_02545_));
 sky130_fd_sc_hd__and3_1 _24471_ (.A(_20313_),
    .B(_20319_),
    .C(_00084_),
    .X(_02689_));
 sky130_vsdinv _24472_ (.A(_19676_),
    .Y(_20320_));
 sky130_fd_sc_hd__buf_2 _24473_ (.A(_20320_),
    .X(_02318_));
 sky130_fd_sc_hd__and3_1 _24474_ (.A(_20318_),
    .B(_02318_),
    .C(_00066_),
    .X(_02544_));
 sky130_fd_sc_hd__and2_1 _24475_ (.A(_02318_),
    .B(_00066_),
    .X(_00067_));
 sky130_fd_sc_hd__and3_1 _24476_ (.A(_00067_),
    .B(_20319_),
    .C(_20313_),
    .X(_02688_));
 sky130_fd_sc_hd__nor2_2 _24477_ (.A(net211),
    .B(net200),
    .Y(_20321_));
 sky130_fd_sc_hd__and3_1 _24478_ (.A(_20318_),
    .B(_20321_),
    .C(_20064_),
    .X(_02543_));
 sky130_vsdinv _24479_ (.A(net306),
    .Y(_20322_));
 sky130_fd_sc_hd__buf_4 _24480_ (.A(_20322_),
    .X(_20323_));
 sky130_fd_sc_hd__nand2_2 _24481_ (.A(_20318_),
    .B(_20321_),
    .Y(_20324_));
 sky130_fd_sc_hd__nor2_1 _24482_ (.A(net226),
    .B(_20324_),
    .Y(_20325_));
 sky130_vsdinv _24483_ (.A(_20325_),
    .Y(_20326_));
 sky130_fd_sc_hd__nor2_1 _24484_ (.A(_20323_),
    .B(_20326_),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_2 _24485_ (.A(\reg_pc[1] ),
    .B(\reg_next_pc[0] ),
    .Y(_20327_));
 sky130_fd_sc_hd__nor2_2 _24486_ (.A(_18525_),
    .B(_20327_),
    .Y(_20328_));
 sky130_fd_sc_hd__and2_1 _24487_ (.A(_20328_),
    .B(net101),
    .X(_20329_));
 sky130_fd_sc_hd__buf_2 _24488_ (.A(_20329_),
    .X(_00307_));
 sky130_fd_sc_hd__and3_1 _24489_ (.A(_18665_),
    .B(_18804_),
    .C(_18595_),
    .X(_00312_));
 sky130_fd_sc_hd__nor2_4 _24490_ (.A(_18532_),
    .B(_18524_),
    .Y(_00303_));
 sky130_vsdinv _24491_ (.A(_00303_),
    .Y(_20330_));
 sky130_fd_sc_hd__nor2_2 _24492_ (.A(_20328_),
    .B(_20330_),
    .Y(_20331_));
 sky130_fd_sc_hd__nor2_2 _24493_ (.A(irq_active),
    .B(\irq_mask[1] ),
    .Y(_20332_));
 sky130_fd_sc_hd__and3_1 _24494_ (.A(_19372_),
    .B(_18677_),
    .C(_20332_),
    .X(_20333_));
 sky130_fd_sc_hd__o211a_1 _24495_ (.A1(_18594_),
    .A2(_00309_),
    .B1(_19597_),
    .C1(_18658_),
    .X(_20334_));
 sky130_fd_sc_hd__a31o_1 _24496_ (.A1(_18541_),
    .A2(_19373_),
    .A3(_20333_),
    .B1(_20334_),
    .X(_20335_));
 sky130_vsdinv _24497_ (.A(\mem_wordsize[2] ),
    .Y(_20336_));
 sky130_fd_sc_hd__nor2_4 _24498_ (.A(_20322_),
    .B(_20336_),
    .Y(_00306_));
 sky130_fd_sc_hd__nor2_2 _24499_ (.A(irq_active),
    .B(\irq_mask[2] ),
    .Y(_20337_));
 sky130_fd_sc_hd__clkbuf_2 _24500_ (.A(_20337_),
    .X(_20338_));
 sky130_vsdinv _24501_ (.A(\mem_wordsize[0] ),
    .Y(_20339_));
 sky130_fd_sc_hd__nor2_8 _24502_ (.A(_20063_),
    .B(_20064_),
    .Y(_00304_));
 sky130_fd_sc_hd__nor2_4 _24503_ (.A(_20339_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__nor2_2 _24504_ (.A(_00306_),
    .B(_00305_),
    .Y(_20340_));
 sky130_fd_sc_hd__o21a_1 _24505_ (.A1(_20340_),
    .A2(_20338_),
    .B1(_03828_),
    .X(_20341_));
 sky130_fd_sc_hd__a31o_1 _24506_ (.A1(_20335_),
    .A2(_00306_),
    .A3(_20338_),
    .B1(_20341_),
    .X(_20342_));
 sky130_fd_sc_hd__nor2_1 _24507_ (.A(_18524_),
    .B(_20340_),
    .Y(_20343_));
 sky130_vsdinv _24508_ (.A(_20337_),
    .Y(_20344_));
 sky130_fd_sc_hd__o21a_1 _24509_ (.A1(_00307_),
    .A2(_20343_),
    .B1(_20344_),
    .X(_20345_));
 sky130_vsdinv _24510_ (.A(_20345_),
    .Y(_20346_));
 sky130_fd_sc_hd__nor2_2 _24511_ (.A(_20330_),
    .B(_20340_),
    .Y(_20347_));
 sky130_fd_sc_hd__o21a_1 _24512_ (.A1(_00307_),
    .A2(_20347_),
    .B1(_20344_),
    .X(_20348_));
 sky130_vsdinv _24513_ (.A(_20348_),
    .Y(_20349_));
 sky130_fd_sc_hd__o211a_1 _24514_ (.A1(_18700_),
    .A2(_18573_),
    .B1(_18768_),
    .C1(_20349_),
    .X(_20350_));
 sky130_vsdinv _24515_ (.A(_20331_),
    .Y(_20351_));
 sky130_fd_sc_hd__nand2_1 _24516_ (.A(_00307_),
    .B(_20344_),
    .Y(_20352_));
 sky130_fd_sc_hd__a311o_1 _24517_ (.A1(_03828_),
    .A2(_20351_),
    .A3(_20352_),
    .B1(_18557_),
    .C1(_00314_),
    .X(_20353_));
 sky130_fd_sc_hd__a311o_1 _24518_ (.A1(_18704_),
    .A2(_18716_),
    .A3(_20346_),
    .B1(_20350_),
    .C1(_20353_),
    .X(_20354_));
 sky130_vsdinv _24519_ (.A(_00306_),
    .Y(_20355_));
 sky130_fd_sc_hd__and2_1 _24520_ (.A(_00305_),
    .B(_20337_),
    .X(_20356_));
 sky130_fd_sc_hd__nand2_1 _24521_ (.A(_20329_),
    .B(_20337_),
    .Y(_20357_));
 sky130_fd_sc_hd__o21ai_1 _24522_ (.A1(_00307_),
    .A2(_20347_),
    .B1(_20357_),
    .Y(_20358_));
 sky130_fd_sc_hd__a31o_1 _24523_ (.A1(_20355_),
    .A2(_20331_),
    .A3(_20356_),
    .B1(_20358_),
    .X(_20359_));
 sky130_fd_sc_hd__a22o_1 _24524_ (.A1(\pcpi_mul.active[1] ),
    .A2(_20349_),
    .B1(_20359_),
    .B2(_20333_),
    .X(_20360_));
 sky130_fd_sc_hd__and3_1 _24525_ (.A(_19373_),
    .B(_18547_),
    .C(_20360_),
    .X(_20361_));
 sky130_fd_sc_hd__nand2_1 _24526_ (.A(_19391_),
    .B(_18594_),
    .Y(_20362_));
 sky130_fd_sc_hd__a21oi_1 _24527_ (.A1(_20362_),
    .A2(_18661_),
    .B1(_20357_),
    .Y(_20363_));
 sky130_fd_sc_hd__a21oi_1 _24528_ (.A1(_00305_),
    .A2(_20344_),
    .B1(_00306_),
    .Y(_20364_));
 sky130_fd_sc_hd__and3_1 _24529_ (.A(_00308_),
    .B(_18540_),
    .C(_20358_),
    .X(_20365_));
 sky130_fd_sc_hd__o31a_1 _24530_ (.A1(_20355_),
    .A2(_20344_),
    .A3(_20330_),
    .B1(_20357_),
    .X(_20366_));
 sky130_fd_sc_hd__or3_4 _24531_ (.A(_00323_),
    .B(_18594_),
    .C(_18662_),
    .X(_20367_));
 sky130_fd_sc_hd__nor2_1 _24532_ (.A(_20366_),
    .B(_20367_),
    .Y(_20368_));
 sky130_fd_sc_hd__a311o_1 _24533_ (.A1(_19393_),
    .A2(_20331_),
    .A3(_20364_),
    .B1(_20365_),
    .C1(_20368_),
    .X(_20369_));
 sky130_vsdinv _24534_ (.A(_20364_),
    .Y(_20370_));
 sky130_fd_sc_hd__a221o_1 _24535_ (.A1(instr_waitirq),
    .A2(do_waitirq),
    .B1(_00303_),
    .B2(_20370_),
    .C1(_20362_),
    .X(_20371_));
 sky130_fd_sc_hd__a21boi_1 _24536_ (.A1(_20355_),
    .A2(_20356_),
    .B1_N(_20343_),
    .Y(_20372_));
 sky130_fd_sc_hd__nand2_1 _24537_ (.A(_20347_),
    .B(_20338_),
    .Y(_20373_));
 sky130_fd_sc_hd__o32a_1 _24538_ (.A1(_18533_),
    .A2(_20372_),
    .A3(_20367_),
    .B1(_18658_),
    .B2(_20373_),
    .X(_20374_));
 sky130_fd_sc_hd__o211a_1 _24539_ (.A1(_19392_),
    .A2(_00303_),
    .B1(_20371_),
    .C1(_20374_),
    .X(_20375_));
 sky130_fd_sc_hd__nor2_1 _24540_ (.A(_00307_),
    .B(_20375_),
    .Y(_20376_));
 sky130_fd_sc_hd__o31a_1 _24541_ (.A1(_20363_),
    .A2(_20369_),
    .A3(_20376_),
    .B1(_19077_),
    .X(_20377_));
 sky130_fd_sc_hd__a2111o_1 _24542_ (.A1(_20331_),
    .A2(_20342_),
    .B1(_20354_),
    .C1(_20361_),
    .D1(_20377_),
    .X(_00039_));
 sky130_fd_sc_hd__nor2_2 _24543_ (.A(_18756_),
    .B(_20345_),
    .Y(_20378_));
 sky130_fd_sc_hd__and2_1 _24544_ (.A(_18784_),
    .B(_20378_),
    .X(_00040_));
 sky130_fd_sc_hd__or2_1 _24545_ (.A(_19360_),
    .B(_18765_),
    .X(_20379_));
 sky130_fd_sc_hd__nand2_1 _24546_ (.A(_18772_),
    .B(_18964_),
    .Y(_20380_));
 sky130_fd_sc_hd__nand2_1 _24547_ (.A(_20380_),
    .B(_18544_),
    .Y(_20381_));
 sky130_vsdinv _24548_ (.A(_20378_),
    .Y(_20382_));
 sky130_fd_sc_hd__a21oi_1 _24549_ (.A1(_20379_),
    .A2(_20381_),
    .B1(_20382_),
    .Y(_00044_));
 sky130_fd_sc_hd__and3_1 _24550_ (.A(_18717_),
    .B(_20306_),
    .C(_01304_),
    .X(_20383_));
 sky130_fd_sc_hd__nand2_1 _24551_ (.A(_18765_),
    .B(_20383_),
    .Y(_20384_));
 sky130_fd_sc_hd__a21oi_1 _24552_ (.A1(_19375_),
    .A2(_20384_),
    .B1(_20382_),
    .Y(_00041_));
 sky130_fd_sc_hd__and4b_1 _24553_ (.A_N(_20332_),
    .B(_19373_),
    .C(_18677_),
    .D(_19372_),
    .X(_20385_));
 sky130_fd_sc_hd__o31a_1 _24554_ (.A1(\cpu_state[0] ),
    .A2(_20345_),
    .A3(_20385_),
    .B1(_19397_),
    .X(_00038_));
 sky130_fd_sc_hd__nand2_1 _24555_ (.A(_20380_),
    .B(\cpu_state[5] ),
    .Y(_20386_));
 sky130_fd_sc_hd__clkbuf_2 _24556_ (.A(_18718_),
    .X(_20387_));
 sky130_fd_sc_hd__buf_4 _24557_ (.A(_20387_),
    .X(_20388_));
 sky130_fd_sc_hd__nand2_1 _24558_ (.A(_19951_),
    .B(_20388_),
    .Y(_20389_));
 sky130_fd_sc_hd__a21oi_1 _24559_ (.A1(_20386_),
    .A2(_20389_),
    .B1(_20382_),
    .Y(_00043_));
 sky130_fd_sc_hd__o21a_4 _24560_ (.A1(mem_do_rdata),
    .A2(_18562_),
    .B1(_18855_),
    .X(net199));
 sky130_vsdinv _24561_ (.A(_19695_),
    .Y(net232));
 sky130_fd_sc_hd__nor2_1 _24562_ (.A(_00291_),
    .B(_20031_),
    .Y(_00317_));
 sky130_fd_sc_hd__clkbuf_4 _24563_ (.A(_18697_),
    .X(_20390_));
 sky130_fd_sc_hd__a32o_1 _24564_ (.A1(_20349_),
    .A2(_18701_),
    .A3(_18773_),
    .B1(alu_wait),
    .B2(_20378_),
    .X(_20391_));
 sky130_fd_sc_hd__a2bb2o_1 _24565_ (.A1_N(_20382_),
    .A2_N(_20308_),
    .B1(_20390_),
    .B2(_20391_),
    .X(_00042_));
 sky130_fd_sc_hd__nor2_2 _24566_ (.A(net200),
    .B(_20322_),
    .Y(_00048_));
 sky130_vsdinv _24567_ (.A(net200),
    .Y(_20392_));
 sky130_fd_sc_hd__nor2_4 _24568_ (.A(net306),
    .B(_20392_),
    .Y(_20393_));
 sky130_fd_sc_hd__nor2_1 _24569_ (.A(_00048_),
    .B(_20393_),
    .Y(_20394_));
 sky130_vsdinv _24570_ (.A(_20394_),
    .Y(_02591_));
 sky130_fd_sc_hd__nor2_1 _24571_ (.A(_19663_),
    .B(net314),
    .Y(_20395_));
 sky130_fd_sc_hd__inv_2 _24572_ (.A(_19663_),
    .Y(_02366_));
 sky130_vsdinv _24573_ (.A(net314),
    .Y(_20396_));
 sky130_fd_sc_hd__nor2_2 _24574_ (.A(_02366_),
    .B(_20396_),
    .Y(_20397_));
 sky130_fd_sc_hd__nor2_2 _24575_ (.A(_20395_),
    .B(_20397_),
    .Y(_20398_));
 sky130_fd_sc_hd__nor2_2 _24576_ (.A(net348),
    .B(_20047_),
    .Y(_20399_));
 sky130_fd_sc_hd__inv_2 _24577_ (.A(net348),
    .Y(_02372_));
 sky130_vsdinv _24578_ (.A(net316),
    .Y(_20400_));
 sky130_fd_sc_hd__nor2_1 _24579_ (.A(_02372_),
    .B(_20400_),
    .Y(_20401_));
 sky130_fd_sc_hd__nor2_2 _24580_ (.A(_20399_),
    .B(_20401_),
    .Y(_20402_));
 sky130_fd_sc_hd__nor2_2 _24581_ (.A(_19662_),
    .B(_20049_),
    .Y(_20403_));
 sky130_fd_sc_hd__inv_2 _24582_ (.A(_19662_),
    .Y(_02369_));
 sky130_vsdinv _24583_ (.A(_20049_),
    .Y(_20404_));
 sky130_fd_sc_hd__nor2_2 _24584_ (.A(_02369_),
    .B(_20404_),
    .Y(_20405_));
 sky130_fd_sc_hd__nor2_2 _24585_ (.A(_20403_),
    .B(_20405_),
    .Y(_20406_));
 sky130_vsdinv _24586_ (.A(_20406_),
    .Y(_20407_));
 sky130_fd_sc_hd__xnor2_1 _24587_ (.A(net345),
    .B(_20050_),
    .Y(_20408_));
 sky130_fd_sc_hd__nand2_1 _24588_ (.A(_20407_),
    .B(_20408_),
    .Y(_20409_));
 sky130_fd_sc_hd__nor2_2 _24589_ (.A(net352),
    .B(_20044_),
    .Y(_20410_));
 sky130_fd_sc_hd__inv_2 _24590_ (.A(net352),
    .Y(_02381_));
 sky130_vsdinv _24591_ (.A(net320),
    .Y(_20411_));
 sky130_fd_sc_hd__nor2_2 _24592_ (.A(_02381_),
    .B(_20411_),
    .Y(_20412_));
 sky130_fd_sc_hd__nor2_2 _24593_ (.A(_20410_),
    .B(_20412_),
    .Y(_20413_));
 sky130_fd_sc_hd__nor2_2 _24594_ (.A(_19660_),
    .B(_20045_),
    .Y(_20414_));
 sky130_fd_sc_hd__inv_2 _24595_ (.A(_19660_),
    .Y(_02378_));
 sky130_vsdinv _24596_ (.A(net319),
    .Y(_20415_));
 sky130_fd_sc_hd__nor2_2 _24597_ (.A(_02378_),
    .B(_20415_),
    .Y(_20416_));
 sky130_fd_sc_hd__nor2_2 _24598_ (.A(_20414_),
    .B(_20416_),
    .Y(_20417_));
 sky130_fd_sc_hd__inv_2 _24599_ (.A(net353),
    .Y(_02384_));
 sky130_vsdinv _24600_ (.A(net321),
    .Y(_20418_));
 sky130_fd_sc_hd__nor2_1 _24601_ (.A(_02384_),
    .B(_20418_),
    .Y(_20419_));
 sky130_vsdinv _24602_ (.A(_20419_),
    .Y(_20420_));
 sky130_fd_sc_hd__nand2_1 _24603_ (.A(_02384_),
    .B(_20418_),
    .Y(_20421_));
 sky130_fd_sc_hd__nand2_1 _24604_ (.A(_20420_),
    .B(_20421_),
    .Y(_20422_));
 sky130_fd_sc_hd__inv_2 _24605_ (.A(net350),
    .Y(_02375_));
 sky130_vsdinv _24606_ (.A(net318),
    .Y(_20423_));
 sky130_fd_sc_hd__nor2_1 _24607_ (.A(_02375_),
    .B(_20423_),
    .Y(_20424_));
 sky130_fd_sc_hd__nand2_1 _24608_ (.A(_02375_),
    .B(_20423_),
    .Y(_20425_));
 sky130_fd_sc_hd__or2b_1 _24609_ (.A(_20424_),
    .B_N(_20425_),
    .X(_20426_));
 sky130_fd_sc_hd__nand2_1 _24610_ (.A(_20422_),
    .B(_20426_),
    .Y(_20427_));
 sky130_fd_sc_hd__or3_1 _24611_ (.A(_20413_),
    .B(_20417_),
    .C(_20427_),
    .X(_20428_));
 sky130_fd_sc_hd__or4_4 _24612_ (.A(_20398_),
    .B(_20402_),
    .C(_20409_),
    .D(_20428_),
    .X(_20429_));
 sky130_fd_sc_hd__nor2_1 _24613_ (.A(_19666_),
    .B(net310),
    .Y(_20430_));
 sky130_fd_sc_hd__inv_2 _24614_ (.A(net342),
    .Y(_02354_));
 sky130_fd_sc_hd__inv_2 _24615_ (.A(net310),
    .Y(_20431_));
 sky130_fd_sc_hd__nor2_1 _24616_ (.A(_02354_),
    .B(_20431_),
    .Y(_20432_));
 sky130_fd_sc_hd__nor2_1 _24617_ (.A(_20430_),
    .B(_20432_),
    .Y(_20433_));
 sky130_vsdinv _24618_ (.A(_20433_),
    .Y(_20434_));
 sky130_fd_sc_hd__nor2_1 _24619_ (.A(net341),
    .B(_20053_),
    .Y(_20435_));
 sky130_fd_sc_hd__inv_2 _24620_ (.A(net341),
    .Y(_02351_));
 sky130_vsdinv _24621_ (.A(net309),
    .Y(_20436_));
 sky130_fd_sc_hd__nor2_1 _24622_ (.A(_02351_),
    .B(_20436_),
    .Y(_20437_));
 sky130_fd_sc_hd__nor2_1 _24623_ (.A(_20435_),
    .B(_20437_),
    .Y(_20438_));
 sky130_vsdinv _24624_ (.A(_20438_),
    .Y(_20439_));
 sky130_fd_sc_hd__nor2_1 _24625_ (.A(net343),
    .B(_20051_),
    .Y(_20440_));
 sky130_fd_sc_hd__inv_2 _24626_ (.A(net343),
    .Y(_02357_));
 sky130_vsdinv _24627_ (.A(net311),
    .Y(_20441_));
 sky130_fd_sc_hd__nor2_1 _24628_ (.A(_02357_),
    .B(_20441_),
    .Y(_20442_));
 sky130_fd_sc_hd__nor2_2 _24629_ (.A(_20440_),
    .B(_20442_),
    .Y(_20443_));
 sky130_vsdinv _24630_ (.A(_20443_),
    .Y(_20444_));
 sky130_fd_sc_hd__inv_2 _24631_ (.A(_19664_),
    .Y(_02360_));
 sky130_fd_sc_hd__clkinv_4 _24632_ (.A(net312),
    .Y(_20445_));
 sky130_fd_sc_hd__nor2_1 _24633_ (.A(_02360_),
    .B(_20445_),
    .Y(_20446_));
 sky130_fd_sc_hd__nand2_1 _24634_ (.A(_02360_),
    .B(_20445_),
    .Y(_20447_));
 sky130_fd_sc_hd__or2b_1 _24635_ (.A(_20446_),
    .B_N(_20447_),
    .X(_20448_));
 sky130_fd_sc_hd__and4_1 _24636_ (.A(_20434_),
    .B(_20439_),
    .C(_20444_),
    .D(_20448_),
    .X(_20449_));
 sky130_vsdinv _24637_ (.A(_20449_),
    .Y(_20450_));
 sky130_fd_sc_hd__nor2_1 _24638_ (.A(_19667_),
    .B(net308),
    .Y(_20451_));
 sky130_fd_sc_hd__inv_2 _24639_ (.A(net340),
    .Y(_02348_));
 sky130_fd_sc_hd__inv_2 _24640_ (.A(net308),
    .Y(_20452_));
 sky130_fd_sc_hd__nor2_1 _24641_ (.A(_02348_),
    .B(_20452_),
    .Y(_20453_));
 sky130_fd_sc_hd__nor2_2 _24642_ (.A(_20451_),
    .B(_20453_),
    .Y(_20454_));
 sky130_fd_sc_hd__nor2_1 _24643_ (.A(_19668_),
    .B(_20055_),
    .Y(_20455_));
 sky130_fd_sc_hd__inv_2 _24644_ (.A(net369),
    .Y(_02342_));
 sky130_vsdinv _24645_ (.A(net337),
    .Y(_20456_));
 sky130_fd_sc_hd__nor2_1 _24646_ (.A(_02342_),
    .B(_20456_),
    .Y(_20457_));
 sky130_fd_sc_hd__nor2_1 _24647_ (.A(_20455_),
    .B(_20457_),
    .Y(_20458_));
 sky130_fd_sc_hd__nor2_1 _24648_ (.A(net368),
    .B(_20056_),
    .Y(_20459_));
 sky130_fd_sc_hd__inv_2 _24649_ (.A(net368),
    .Y(_02339_));
 sky130_vsdinv _24650_ (.A(net336),
    .Y(_20460_));
 sky130_fd_sc_hd__nor2_1 _24651_ (.A(_02339_),
    .B(_20460_),
    .Y(_20461_));
 sky130_fd_sc_hd__nor2_1 _24652_ (.A(_20459_),
    .B(_20461_),
    .Y(_20462_));
 sky130_fd_sc_hd__nor2_1 _24653_ (.A(net339),
    .B(_20054_),
    .Y(_20463_));
 sky130_fd_sc_hd__inv_2 _24654_ (.A(net339),
    .Y(_02345_));
 sky130_vsdinv _24655_ (.A(net307),
    .Y(_20464_));
 sky130_fd_sc_hd__nor2_2 _24656_ (.A(_02345_),
    .B(_20464_),
    .Y(_20465_));
 sky130_fd_sc_hd__nor2_2 _24657_ (.A(_20463_),
    .B(_20465_),
    .Y(_20466_));
 sky130_fd_sc_hd__or4_4 _24658_ (.A(_20454_),
    .B(_20458_),
    .C(_20462_),
    .D(_20466_),
    .X(_20467_));
 sky130_fd_sc_hd__nor2_2 _24659_ (.A(net227),
    .B(_20059_),
    .Y(_20468_));
 sky130_fd_sc_hd__inv_2 _24660_ (.A(net227),
    .Y(_02330_));
 sky130_vsdinv _24661_ (.A(net333),
    .Y(_20469_));
 sky130_fd_sc_hd__nor2_2 _24662_ (.A(_02330_),
    .B(_20469_),
    .Y(_20470_));
 sky130_fd_sc_hd__nor2_2 _24663_ (.A(_20468_),
    .B(_20470_),
    .Y(_20471_));
 sky130_fd_sc_hd__inv_2 _24664_ (.A(net228),
    .Y(_02333_));
 sky130_vsdinv _24665_ (.A(net334),
    .Y(_20472_));
 sky130_fd_sc_hd__nor2_1 _24666_ (.A(_02333_),
    .B(_20472_),
    .Y(_20473_));
 sky130_fd_sc_hd__nand2_1 _24667_ (.A(_02333_),
    .B(_20472_),
    .Y(_20474_));
 sky130_fd_sc_hd__or2b_1 _24668_ (.A(_20473_),
    .B_N(_20474_),
    .X(_20475_));
 sky130_vsdinv _24669_ (.A(_20475_),
    .Y(_20476_));
 sky130_fd_sc_hd__nor2_1 _24670_ (.A(net225),
    .B(_20061_),
    .Y(_20477_));
 sky130_fd_sc_hd__inv_2 _24671_ (.A(net225),
    .Y(_02324_));
 sky130_vsdinv _24672_ (.A(_20061_),
    .Y(_20478_));
 sky130_fd_sc_hd__nor2_2 _24673_ (.A(_02324_),
    .B(_20478_),
    .Y(_20479_));
 sky130_fd_sc_hd__nor2_2 _24674_ (.A(_20477_),
    .B(_20479_),
    .Y(_20480_));
 sky130_fd_sc_hd__nor2_1 _24675_ (.A(net222),
    .B(_20062_),
    .Y(_20481_));
 sky130_vsdinv _24676_ (.A(net328),
    .Y(_20482_));
 sky130_fd_sc_hd__nor2_1 _24677_ (.A(_20319_),
    .B(_20482_),
    .Y(_20483_));
 sky130_fd_sc_hd__nor2_1 _24678_ (.A(_20481_),
    .B(_20483_),
    .Y(_20484_));
 sky130_fd_sc_hd__nor2_1 _24679_ (.A(_20480_),
    .B(_20484_),
    .Y(_20485_));
 sky130_fd_sc_hd__or3b_1 _24680_ (.A(_20471_),
    .B(_20476_),
    .C_N(_20485_),
    .X(_20486_));
 sky130_fd_sc_hd__nor2_1 _24681_ (.A(net226),
    .B(_20060_),
    .Y(_20487_));
 sky130_vsdinv _24682_ (.A(net332),
    .Y(_20488_));
 sky130_fd_sc_hd__nor2_1 _24683_ (.A(_20309_),
    .B(_20488_),
    .Y(_20489_));
 sky130_fd_sc_hd__nor2_1 _24684_ (.A(_20487_),
    .B(_20489_),
    .Y(_20490_));
 sky130_vsdinv _24685_ (.A(_20490_),
    .Y(_20491_));
 sky130_vsdinv _24686_ (.A(_20063_),
    .Y(_20492_));
 sky130_fd_sc_hd__nor2_1 _24687_ (.A(_20320_),
    .B(_20492_),
    .Y(_20493_));
 sky130_fd_sc_hd__buf_6 _24688_ (.A(_20492_),
    .X(_20494_));
 sky130_fd_sc_hd__nand2_1 _24689_ (.A(_02318_),
    .B(_20494_),
    .Y(_20495_));
 sky130_fd_sc_hd__or2b_1 _24690_ (.A(_20493_),
    .B_N(_20495_),
    .X(_20496_));
 sky130_fd_sc_hd__xnor2_1 _24691_ (.A(net229),
    .B(_20057_),
    .Y(_20497_));
 sky130_fd_sc_hd__and4_1 _24692_ (.A(_20491_),
    .B(_20394_),
    .C(_20496_),
    .D(_20497_),
    .X(_20498_));
 sky130_fd_sc_hd__or4b_4 _24693_ (.A(_20450_),
    .B(_20467_),
    .C(_20486_),
    .D_N(_20498_),
    .X(_20499_));
 sky130_fd_sc_hd__nor2_1 _24694_ (.A(_19659_),
    .B(_20040_),
    .Y(_20500_));
 sky130_fd_sc_hd__inv_2 _24695_ (.A(net355),
    .Y(_02390_));
 sky130_vsdinv _24696_ (.A(net323),
    .Y(_20501_));
 sky130_fd_sc_hd__nor2_1 _24697_ (.A(_02390_),
    .B(_20501_),
    .Y(_20502_));
 sky130_fd_sc_hd__nor2_2 _24698_ (.A(_20500_),
    .B(_20502_),
    .Y(_20503_));
 sky130_fd_sc_hd__nor2_1 _24699_ (.A(net358),
    .B(_20038_),
    .Y(_20504_));
 sky130_fd_sc_hd__inv_2 _24700_ (.A(net358),
    .Y(_02399_));
 sky130_fd_sc_hd__clkinv_4 _24701_ (.A(net326),
    .Y(_20505_));
 sky130_fd_sc_hd__nor2_1 _24702_ (.A(_02399_),
    .B(_20505_),
    .Y(_20506_));
 sky130_fd_sc_hd__nor2_2 _24703_ (.A(_20504_),
    .B(_20506_),
    .Y(_20507_));
 sky130_fd_sc_hd__nor2_1 _24704_ (.A(_19657_),
    .B(_20039_),
    .Y(_20508_));
 sky130_fd_sc_hd__inv_2 _24705_ (.A(net356),
    .Y(_02393_));
 sky130_vsdinv _24706_ (.A(net324),
    .Y(_20509_));
 sky130_fd_sc_hd__nor2_1 _24707_ (.A(_02393_),
    .B(_20509_),
    .Y(_20510_));
 sky130_fd_sc_hd__nor2_2 _24708_ (.A(_20508_),
    .B(_20510_),
    .Y(_20511_));
 sky130_fd_sc_hd__nor2_1 _24709_ (.A(net354),
    .B(_20042_),
    .Y(_20512_));
 sky130_fd_sc_hd__inv_2 _24710_ (.A(net354),
    .Y(_02387_));
 sky130_vsdinv _24711_ (.A(_20042_),
    .Y(_20513_));
 sky130_fd_sc_hd__nor2_1 _24712_ (.A(_02387_),
    .B(_20513_),
    .Y(_20514_));
 sky130_fd_sc_hd__nor2_1 _24713_ (.A(_20512_),
    .B(_20514_),
    .Y(_20515_));
 sky130_fd_sc_hd__or4_4 _24714_ (.A(_20503_),
    .B(_20507_),
    .C(_20511_),
    .D(_20515_),
    .X(_20516_));
 sky130_fd_sc_hd__nor2_1 _24715_ (.A(_19655_),
    .B(net327),
    .Y(_20517_));
 sky130_fd_sc_hd__inv_2 _24716_ (.A(net359),
    .Y(_02402_));
 sky130_vsdinv _24717_ (.A(net327),
    .Y(_20518_));
 sky130_fd_sc_hd__nor2_2 _24718_ (.A(_02402_),
    .B(_20518_),
    .Y(_20519_));
 sky130_fd_sc_hd__nor2_2 _24719_ (.A(_20517_),
    .B(_20519_),
    .Y(_20520_));
 sky130_fd_sc_hd__nor2_1 _24720_ (.A(_19656_),
    .B(net325),
    .Y(_20521_));
 sky130_fd_sc_hd__inv_2 _24721_ (.A(net357),
    .Y(_02396_));
 sky130_vsdinv _24722_ (.A(net325),
    .Y(_20522_));
 sky130_fd_sc_hd__nor2_1 _24723_ (.A(_02396_),
    .B(_20522_),
    .Y(_20523_));
 sky130_fd_sc_hd__nor2_2 _24724_ (.A(_20521_),
    .B(_20523_),
    .Y(_20524_));
 sky130_fd_sc_hd__nor2_2 _24725_ (.A(net330),
    .B(net362),
    .Y(_20525_));
 sky130_fd_sc_hd__nor2_4 _24726_ (.A(_18667_),
    .B(_18690_),
    .Y(_20526_));
 sky130_fd_sc_hd__nor2_4 _24727_ (.A(_20525_),
    .B(_20526_),
    .Y(_20527_));
 sky130_fd_sc_hd__nor2_2 _24728_ (.A(net361),
    .B(_20036_),
    .Y(_20528_));
 sky130_fd_sc_hd__inv_2 _24729_ (.A(net361),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _24730_ (.A(net329),
    .Y(_20529_));
 sky130_fd_sc_hd__nor2_2 _24731_ (.A(_02405_),
    .B(_20529_),
    .Y(_20530_));
 sky130_fd_sc_hd__nor2_2 _24732_ (.A(_20528_),
    .B(_20530_),
    .Y(_20531_));
 sky130_fd_sc_hd__or4_4 _24733_ (.A(_20520_),
    .B(_20524_),
    .C(_20527_),
    .D(_20531_),
    .X(_20532_));
 sky130_fd_sc_hd__nor2_1 _24734_ (.A(_20516_),
    .B(_20532_),
    .Y(_20533_));
 sky130_fd_sc_hd__nor3b_4 _24735_ (.A(_20429_),
    .B(_20499_),
    .C_N(_20533_),
    .Y(_00000_));
 sky130_fd_sc_hd__and3_1 _24736_ (.A(_18672_),
    .B(_18675_),
    .C(_18683_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_1 _24737_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00006_));
 sky130_fd_sc_hd__or3_1 _24738_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00007_));
 sky130_fd_sc_hd__nand2_1 _24739_ (.A(_18569_),
    .B(_20193_),
    .Y(_00299_));
 sky130_fd_sc_hd__a2111o_1 _24740_ (.A1(_18721_),
    .A2(_00297_),
    .B1(_18533_),
    .C1(_00319_),
    .D1(_00317_),
    .X(_20534_));
 sky130_fd_sc_hd__a31oi_2 _24741_ (.A1(mem_do_prefetch),
    .A2(_18530_),
    .A3(_18777_),
    .B1(_20534_),
    .Y(_20535_));
 sky130_fd_sc_hd__nor2_1 _24742_ (.A(_18853_),
    .B(_18756_),
    .Y(_20536_));
 sky130_fd_sc_hd__or2_1 _24743_ (.A(instr_lhu),
    .B(instr_lh),
    .X(_20537_));
 sky130_fd_sc_hd__a32o_1 _24744_ (.A1(instr_sh),
    .A2(\cpu_state[5] ),
    .A3(_20536_),
    .B1(_18966_),
    .B2(_20537_),
    .X(_20538_));
 sky130_fd_sc_hd__a2bb2o_1 _24745_ (.A1_N(_20336_),
    .A2_N(_20535_),
    .B1(_18965_),
    .B2(_20538_),
    .X(_00047_));
 sky130_fd_sc_hd__clkbuf_4 _24746_ (.A(_18767_),
    .X(_20539_));
 sky130_fd_sc_hd__clkbuf_4 _24747_ (.A(_20539_),
    .X(_20540_));
 sky130_fd_sc_hd__buf_4 _24748_ (.A(_18960_),
    .X(_20541_));
 sky130_fd_sc_hd__and3_1 _24749_ (.A(_20540_),
    .B(_20541_),
    .C(_20031_),
    .X(_00336_));
 sky130_fd_sc_hd__o21ai_1 _24750_ (.A1(mem_do_rinst),
    .A2(_18964_),
    .B1(_18573_),
    .Y(_00338_));
 sky130_vsdinv _24751_ (.A(alu_eq),
    .Y(_00340_));
 sky130_fd_sc_hd__or3_4 _24752_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .C(is_sltiu_bltu_sltu),
    .X(_20542_));
 sky130_fd_sc_hd__nor3_4 _24753_ (.A(instr_bgeu),
    .B(instr_bge),
    .C(_20542_),
    .Y(_00341_));
 sky130_vsdinv _24754_ (.A(instr_bge),
    .Y(_20543_));
 sky130_fd_sc_hd__nand2_1 _24755_ (.A(is_sltiu_bltu_sltu),
    .B(alu_ltu),
    .Y(_20544_));
 sky130_fd_sc_hd__nand2_1 _24756_ (.A(is_slti_blt_slt),
    .B(alu_lts),
    .Y(_20545_));
 sky130_fd_sc_hd__o221a_1 _24757_ (.A1(alu_eq),
    .A2(_18948_),
    .B1(_18941_),
    .B2(alu_ltu),
    .C1(_20545_),
    .X(_20546_));
 sky130_fd_sc_hd__o211a_1 _24758_ (.A1(_20543_),
    .A2(alu_lts),
    .B1(_20544_),
    .C1(_20546_),
    .X(_00342_));
 sky130_fd_sc_hd__nand2_1 _24759_ (.A(_21108_),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__o22ai_1 _24760_ (.A1(_00346_),
    .A2(_20540_),
    .B1(_00339_),
    .B2(_00297_),
    .Y(_00347_));
 sky130_fd_sc_hd__nor2_1 _24761_ (.A(_18761_),
    .B(_18660_),
    .Y(_00349_));
 sky130_fd_sc_hd__and2_1 _24762_ (.A(_02410_),
    .B(_00349_),
    .X(_00351_));
 sky130_fd_sc_hd__o21a_1 _24763_ (.A1(_20540_),
    .A2(_18964_),
    .B1(_18959_),
    .X(_00355_));
 sky130_fd_sc_hd__inv_2 _24764_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_vsdinv _24765_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_vsdinv _24766_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_vsdinv _24767_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_vsdinv _24768_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_vsdinv _24769_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_vsdinv _24770_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_vsdinv _24771_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_vsdinv _24772_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_vsdinv _24773_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_vsdinv _24774_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_vsdinv _24775_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_vsdinv _24776_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_vsdinv _24777_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_vsdinv _24778_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_vsdinv _24779_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_vsdinv _24780_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_vsdinv _24781_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_vsdinv _24782_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_vsdinv _24783_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_vsdinv _24784_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_vsdinv _24785_ (.A(alu_wait),
    .Y(_00302_));
 sky130_vsdinv _24786_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_vsdinv _24787_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_vsdinv _24788_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_vsdinv _24789_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_vsdinv _24790_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_vsdinv _24791_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_vsdinv _24792_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_vsdinv _24793_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_vsdinv _24794_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_vsdinv _24795_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_vsdinv _24796_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_vsdinv _24797_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_vsdinv _24798_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_vsdinv _24799_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_vsdinv _24800_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_vsdinv _24801_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_vsdinv _24802_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_vsdinv _24803_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_vsdinv _24804_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_vsdinv _24805_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_vsdinv _24806_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_vsdinv _24807_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_vsdinv _24808_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_vsdinv _24809_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_vsdinv _24810_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_vsdinv _24811_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_vsdinv _24812_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_vsdinv _24813_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_vsdinv _24814_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_vsdinv _24815_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_vsdinv _24816_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_vsdinv _24817_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_vsdinv _24818_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_vsdinv _24819_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_vsdinv _24820_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_vsdinv _24821_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_vsdinv _24822_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_vsdinv _24823_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_vsdinv _24824_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_vsdinv _24825_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_vsdinv _24826_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_vsdinv _24827_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_vsdinv _24828_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_vsdinv _24829_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_vsdinv _24830_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_vsdinv _24831_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_vsdinv _24832_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_vsdinv _24833_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_vsdinv _24834_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_vsdinv _24835_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_vsdinv _24836_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_vsdinv _24837_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_vsdinv _24838_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_vsdinv _24839_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_vsdinv _24840_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_vsdinv _24841_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_vsdinv _24842_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_vsdinv _24843_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_vsdinv _24844_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_vsdinv _24845_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_vsdinv _24846_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_vsdinv _24847_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_vsdinv _24848_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_vsdinv _24849_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_vsdinv _24850_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_vsdinv _24851_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_vsdinv _24852_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_vsdinv _24853_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_vsdinv _24854_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_vsdinv _24855_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_vsdinv _24856_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_vsdinv _24857_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_vsdinv _24858_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_vsdinv _24859_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_vsdinv _24860_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_vsdinv _24861_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_vsdinv _24862_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_vsdinv _24863_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_vsdinv _24864_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_vsdinv _24865_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_vsdinv _24866_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_vsdinv _24867_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_vsdinv _24868_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_vsdinv _24869_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_vsdinv _24870_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_vsdinv _24871_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_vsdinv _24872_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_vsdinv _24873_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_vsdinv _24874_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_vsdinv _24875_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_vsdinv _24876_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_vsdinv _24877_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_vsdinv _24878_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_vsdinv _24879_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_vsdinv _24880_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_vsdinv _24881_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_vsdinv _24882_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_vsdinv _24883_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_vsdinv _24884_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_vsdinv _24885_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_vsdinv _24886_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_vsdinv _24887_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_vsdinv _24888_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_vsdinv _24889_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_vsdinv _24890_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_vsdinv _24891_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_vsdinv _24892_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_vsdinv _24893_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_vsdinv _24894_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_vsdinv _24895_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_vsdinv _24896_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_vsdinv _24897_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_vsdinv _24898_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_vsdinv _24899_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_vsdinv _24900_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_vsdinv _24901_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_vsdinv _24902_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_vsdinv _24903_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_vsdinv _24904_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_vsdinv _24905_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_vsdinv _24906_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_vsdinv _24907_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_vsdinv _24908_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_vsdinv _24909_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_vsdinv _24910_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_vsdinv _24911_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_vsdinv _24912_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_vsdinv _24913_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_vsdinv _24914_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_vsdinv _24915_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_vsdinv _24916_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_vsdinv _24917_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_vsdinv _24918_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_vsdinv _24919_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_vsdinv _24920_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_vsdinv _24921_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_vsdinv _24922_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_vsdinv _24923_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_vsdinv _24924_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_vsdinv _24925_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_vsdinv _24926_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_vsdinv _24927_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_vsdinv _24928_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_vsdinv _24929_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_vsdinv _24930_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_vsdinv _24931_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_vsdinv _24932_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_vsdinv _24933_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_vsdinv _24934_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_vsdinv _24935_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_vsdinv _24936_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_vsdinv _24937_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_vsdinv _24938_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_vsdinv _24939_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_vsdinv _24940_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_vsdinv _24941_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_vsdinv _24942_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_vsdinv _24943_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_vsdinv _24944_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_vsdinv _24945_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_vsdinv _24946_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_vsdinv _24947_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_vsdinv _24948_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_vsdinv _24949_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_vsdinv _24950_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_vsdinv _24951_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_vsdinv _24952_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_vsdinv _24953_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_vsdinv _24954_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_vsdinv _24955_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_vsdinv _24956_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_vsdinv _24957_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_vsdinv _24958_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_vsdinv _24959_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_vsdinv _24960_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_vsdinv _24961_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_vsdinv _24962_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_vsdinv _24963_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_vsdinv _24964_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_vsdinv _24965_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_vsdinv _24966_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_vsdinv _24967_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_vsdinv _24968_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_vsdinv _24969_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_vsdinv _24970_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_vsdinv _24971_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_vsdinv _24972_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_vsdinv _24973_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_vsdinv _24974_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_vsdinv _24975_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_vsdinv _24976_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_vsdinv _24977_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_vsdinv _24978_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_vsdinv _24979_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_vsdinv _24980_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_vsdinv _24981_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_vsdinv _24982_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_vsdinv _24983_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_vsdinv _24984_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_vsdinv _24985_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_vsdinv _24986_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_vsdinv _24987_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_vsdinv _24988_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_vsdinv _24989_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_vsdinv _24990_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_vsdinv _24991_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_vsdinv _24992_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_vsdinv _24993_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_vsdinv _24994_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_vsdinv _24995_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_vsdinv _24996_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_vsdinv _24997_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_vsdinv _24998_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_vsdinv _24999_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_vsdinv _25000_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_vsdinv _25001_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_vsdinv _25002_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_vsdinv _25003_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_vsdinv _25004_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_vsdinv _25005_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_vsdinv _25006_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_vsdinv _25007_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_vsdinv _25008_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_vsdinv _25009_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_vsdinv _25010_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_vsdinv _25011_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_vsdinv _25012_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_vsdinv _25013_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_vsdinv _25014_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_vsdinv _25015_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_vsdinv _25016_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_vsdinv _25017_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_vsdinv _25018_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_vsdinv _25019_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_vsdinv _25020_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_vsdinv _25021_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_vsdinv _25022_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_vsdinv _25023_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_vsdinv _25024_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_vsdinv _25025_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_vsdinv _25026_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_vsdinv _25027_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_vsdinv _25028_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_vsdinv _25029_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_vsdinv _25030_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_vsdinv _25031_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_vsdinv _25032_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_vsdinv _25033_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_vsdinv _25034_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_vsdinv _25035_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_vsdinv _25036_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_vsdinv _25037_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_vsdinv _25038_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_vsdinv _25039_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_vsdinv _25040_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_vsdinv _25041_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_vsdinv _25042_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_vsdinv _25043_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_vsdinv _25044_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_vsdinv _25045_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_vsdinv _25046_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_vsdinv _25047_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_vsdinv _25048_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_vsdinv _25049_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_vsdinv _25050_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_vsdinv _25051_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_vsdinv _25052_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_vsdinv _25053_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_vsdinv _25054_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_vsdinv _25055_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_vsdinv _25056_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_vsdinv _25057_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_vsdinv _25058_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_vsdinv _25059_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_vsdinv _25060_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_vsdinv _25061_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_vsdinv _25062_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_vsdinv _25063_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_vsdinv _25064_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_vsdinv _25065_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_vsdinv _25066_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_vsdinv _25067_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_vsdinv _25068_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_vsdinv _25069_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_vsdinv _25070_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_vsdinv _25071_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_vsdinv _25072_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_vsdinv _25073_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_vsdinv _25074_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_vsdinv _25075_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_vsdinv _25076_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_vsdinv _25077_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_vsdinv _25078_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_vsdinv _25079_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_vsdinv _25080_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_vsdinv _25081_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_vsdinv _25082_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_vsdinv _25083_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_vsdinv _25084_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_vsdinv _25085_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_vsdinv _25086_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_vsdinv _25087_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_vsdinv _25088_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_vsdinv _25089_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_vsdinv _25090_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_vsdinv _25091_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_vsdinv _25092_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_vsdinv _25093_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_vsdinv _25094_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_vsdinv _25095_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_vsdinv _25096_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_vsdinv _25097_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_vsdinv _25098_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_vsdinv _25099_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_vsdinv _25100_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_vsdinv _25101_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_vsdinv _25102_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_vsdinv _25103_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_vsdinv _25104_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_vsdinv _25105_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_vsdinv _25106_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_vsdinv _25107_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_vsdinv _25108_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_vsdinv _25109_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_vsdinv _25110_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_vsdinv _25111_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_vsdinv _25112_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_vsdinv _25113_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_vsdinv _25114_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_vsdinv _25115_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_vsdinv _25116_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_vsdinv _25117_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_vsdinv _25118_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_vsdinv _25119_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_vsdinv _25120_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_vsdinv _25121_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_vsdinv _25122_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_vsdinv _25123_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_vsdinv _25124_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_vsdinv _25125_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_vsdinv _25126_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_vsdinv _25127_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_vsdinv _25128_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_vsdinv _25129_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_vsdinv _25130_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_vsdinv _25131_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_vsdinv _25132_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_vsdinv _25133_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_vsdinv _25134_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_vsdinv _25135_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_vsdinv _25136_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_vsdinv _25137_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_vsdinv _25138_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_vsdinv _25139_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_vsdinv _25140_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_vsdinv _25141_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_vsdinv _25142_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_vsdinv _25143_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_vsdinv _25144_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_vsdinv _25145_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_vsdinv _25146_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_vsdinv _25147_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_vsdinv _25148_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_vsdinv _25149_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_vsdinv _25150_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_vsdinv _25151_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_vsdinv _25152_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_vsdinv _25153_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_vsdinv _25154_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_vsdinv _25155_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_vsdinv _25156_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_vsdinv _25157_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_vsdinv _25158_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_vsdinv _25159_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_vsdinv _25160_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_vsdinv _25161_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_vsdinv _25162_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_vsdinv _25163_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_vsdinv _25164_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_vsdinv _25165_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_vsdinv _25166_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_vsdinv _25167_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_vsdinv _25168_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_vsdinv _25169_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_vsdinv _25170_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_vsdinv _25171_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_vsdinv _25172_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_vsdinv _25173_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_vsdinv _25174_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_vsdinv _25175_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_vsdinv _25176_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_vsdinv _25177_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_vsdinv _25178_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_vsdinv _25179_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_vsdinv _25180_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_vsdinv _25181_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_vsdinv _25182_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_vsdinv _25183_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_vsdinv _25184_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_vsdinv _25185_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_vsdinv _25186_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_vsdinv _25187_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_vsdinv _25188_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_vsdinv _25189_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_vsdinv _25190_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_vsdinv _25191_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_vsdinv _25192_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_vsdinv _25193_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__a32o_1 _25194_ (.A1(instr_sw),
    .A2(\cpu_state[5] ),
    .A3(_20536_),
    .B1(_18966_),
    .B2(instr_lw),
    .X(_20547_));
 sky130_fd_sc_hd__nor2_1 _25195_ (.A(_20339_),
    .B(_20535_),
    .Y(_20548_));
 sky130_fd_sc_hd__a211o_1 _25196_ (.A1(_18965_),
    .A2(_20547_),
    .B1(_19597_),
    .C1(_20548_),
    .X(_00045_));
 sky130_vsdinv _25197_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_vsdinv _25198_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_vsdinv _25199_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_vsdinv _25200_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_vsdinv _25201_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_vsdinv _25202_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_vsdinv _25203_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_vsdinv _25204_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_vsdinv _25205_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_vsdinv _25206_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_vsdinv _25207_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_vsdinv _25208_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_vsdinv _25209_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_vsdinv _25210_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_vsdinv _25211_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_vsdinv _25212_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_vsdinv _25213_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_vsdinv _25214_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_vsdinv _25215_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_vsdinv _25216_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_vsdinv _25217_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_vsdinv _25218_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_vsdinv _25219_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_vsdinv _25220_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_vsdinv _25221_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_vsdinv _25222_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_vsdinv _25223_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_vsdinv _25224_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_vsdinv _25225_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_vsdinv _25226_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_vsdinv _25227_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_vsdinv _25228_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_vsdinv _25229_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_vsdinv _25230_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_vsdinv _25231_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_vsdinv _25232_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_vsdinv _25233_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_vsdinv _25234_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_vsdinv _25235_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_vsdinv _25236_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_vsdinv _25237_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_vsdinv _25238_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_vsdinv _25239_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_vsdinv _25240_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_vsdinv _25241_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_vsdinv _25242_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_vsdinv _25243_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_vsdinv _25244_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_vsdinv _25245_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_vsdinv _25246_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_vsdinv _25247_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_vsdinv _25248_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_vsdinv _25249_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_vsdinv _25250_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_vsdinv _25251_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_vsdinv _25252_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_vsdinv _25253_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_vsdinv _25254_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_vsdinv _25255_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_vsdinv _25256_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2_2 _25257_ (.A(\mem_state[1] ),
    .B(_18571_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _25258_ (.A(_18569_),
    .B(_00289_),
    .Y(_00298_));
 sky130_vsdinv _25259_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_vsdinv _25260_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_vsdinv _25261_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_vsdinv _25262_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_vsdinv _25263_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_vsdinv _25264_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_vsdinv _25265_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_vsdinv _25266_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_vsdinv _25267_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_vsdinv _25268_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_vsdinv _25269_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_vsdinv _25270_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_vsdinv _25271_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_vsdinv _25272_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_vsdinv _25273_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_vsdinv _25274_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_vsdinv _25275_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_vsdinv _25276_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_vsdinv _25277_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_vsdinv _25278_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_vsdinv _25279_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_vsdinv _25280_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_vsdinv _25281_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_vsdinv _25282_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_vsdinv _25283_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_vsdinv _25284_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_vsdinv _25285_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_vsdinv _25286_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_vsdinv _25287_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_vsdinv _25288_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_vsdinv _25289_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_vsdinv _25290_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_vsdinv _25291_ (.A(\mem_wordsize[1] ),
    .Y(_20549_));
 sky130_fd_sc_hd__clkbuf_2 _25292_ (.A(_20549_),
    .X(_20550_));
 sky130_fd_sc_hd__clkbuf_2 _25293_ (.A(_18535_),
    .X(_20551_));
 sky130_fd_sc_hd__o211a_1 _25294_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_18544_),
    .C1(_20551_),
    .X(_20552_));
 sky130_fd_sc_hd__a31o_1 _25295_ (.A1(_00291_),
    .A2(instr_sb),
    .A3(\cpu_state[5] ),
    .B1(_20552_),
    .X(_20553_));
 sky130_fd_sc_hd__a2bb2o_1 _25296_ (.A1_N(_20550_),
    .A2_N(_20535_),
    .B1(_18534_),
    .B2(_20553_),
    .X(_00046_));
 sky130_vsdinv _25297_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_vsdinv _25298_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_vsdinv _25299_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_vsdinv _25300_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_vsdinv _25301_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_vsdinv _25302_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_vsdinv _25303_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_vsdinv _25304_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_vsdinv _25305_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_vsdinv _25306_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_vsdinv _25307_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_vsdinv _25308_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_vsdinv _25309_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_vsdinv _25310_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_vsdinv _25311_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_vsdinv _25312_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_vsdinv _25313_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_vsdinv _25314_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_vsdinv _25315_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_vsdinv _25316_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_vsdinv _25317_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_vsdinv _25318_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_vsdinv _25319_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_vsdinv _25320_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_vsdinv _25321_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_vsdinv _25322_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_vsdinv _25323_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_vsdinv _25324_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_vsdinv _25325_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_vsdinv _25326_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_vsdinv _25327_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_vsdinv _25328_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_vsdinv _25329_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_vsdinv _25330_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_vsdinv _25331_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_vsdinv _25332_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_vsdinv _25333_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_vsdinv _25334_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_vsdinv _25335_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_vsdinv _25336_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_vsdinv _25337_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_vsdinv _25338_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_vsdinv _25339_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_vsdinv _25340_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_vsdinv _25341_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_vsdinv _25342_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_vsdinv _25343_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_vsdinv _25344_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_vsdinv _25345_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_vsdinv _25346_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_vsdinv _25347_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_vsdinv _25348_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_vsdinv _25349_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_vsdinv _25350_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__clkbuf_4 _25351_ (.A(latched_branch),
    .X(_20554_));
 sky130_fd_sc_hd__clkbuf_4 _25352_ (.A(_20554_),
    .X(_20555_));
 sky130_fd_sc_hd__and2_1 _25353_ (.A(_20555_),
    .B(_00294_),
    .X(_00295_));
 sky130_vsdinv _25354_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_vsdinv _25355_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_vsdinv _25356_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_vsdinv _25357_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_vsdinv _25358_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_vsdinv _25359_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_vsdinv _25360_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_vsdinv _25361_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_vsdinv _25362_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_vsdinv _25363_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_vsdinv _25364_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_vsdinv _25365_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_vsdinv _25366_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_vsdinv _25367_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_vsdinv _25368_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_vsdinv _25369_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_vsdinv _25370_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_vsdinv _25371_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_vsdinv _25372_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_vsdinv _25373_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_vsdinv _25374_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_vsdinv _25375_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_vsdinv _25376_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_vsdinv _25377_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_vsdinv _25378_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_vsdinv _25379_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_vsdinv _25380_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_vsdinv _25381_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_vsdinv _25382_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_vsdinv _25383_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_vsdinv _25384_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_vsdinv _25385_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_vsdinv _25386_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_vsdinv _25387_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_vsdinv _25388_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_vsdinv _25389_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_vsdinv _25390_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_vsdinv _25391_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_vsdinv _25392_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_vsdinv _25393_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_vsdinv _25394_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_vsdinv _25395_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_vsdinv _25396_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_vsdinv _25397_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_vsdinv _25398_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_vsdinv _25399_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_fd_sc_hd__or4_4 _25400_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_20556_));
 sky130_fd_sc_hd__nor2_1 _25401_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .Y(_20557_));
 sky130_vsdinv _25402_ (.A(_20557_),
    .Y(_20558_));
 sky130_fd_sc_hd__or2_1 _25403_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .X(_20559_));
 sky130_fd_sc_hd__nor2_1 _25404_ (.A(\timer[2] ),
    .B(_20559_),
    .Y(_20560_));
 sky130_vsdinv _25405_ (.A(\timer[3] ),
    .Y(_20561_));
 sky130_fd_sc_hd__nand2_1 _25406_ (.A(_20560_),
    .B(_20561_),
    .Y(_20562_));
 sky130_fd_sc_hd__nor2_1 _25407_ (.A(_20558_),
    .B(_20562_),
    .Y(_20563_));
 sky130_vsdinv _25408_ (.A(_20563_),
    .Y(_20564_));
 sky130_fd_sc_hd__nor2_1 _25409_ (.A(\timer[6] ),
    .B(_20564_),
    .Y(_20565_));
 sky130_vsdinv _25410_ (.A(_20565_),
    .Y(_20566_));
 sky130_fd_sc_hd__nor2_2 _25411_ (.A(\timer[7] ),
    .B(_20566_),
    .Y(_20567_));
 sky130_fd_sc_hd__nor2_1 _25412_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .Y(_20568_));
 sky130_fd_sc_hd__nand2_1 _25413_ (.A(_20567_),
    .B(_20568_),
    .Y(_20569_));
 sky130_fd_sc_hd__or2_1 _25414_ (.A(\timer[10] ),
    .B(_20569_),
    .X(_20570_));
 sky130_fd_sc_hd__or2_1 _25415_ (.A(\timer[11] ),
    .B(_20570_),
    .X(_20571_));
 sky130_fd_sc_hd__or2_1 _25416_ (.A(\timer[12] ),
    .B(_20571_),
    .X(_20572_));
 sky130_fd_sc_hd__nor2_2 _25417_ (.A(\timer[13] ),
    .B(_20572_),
    .Y(_20573_));
 sky130_vsdinv _25418_ (.A(\timer[14] ),
    .Y(_20574_));
 sky130_fd_sc_hd__nand2_2 _25419_ (.A(_20573_),
    .B(_20574_),
    .Y(_20575_));
 sky130_fd_sc_hd__nor2_4 _25420_ (.A(\timer[15] ),
    .B(_20575_),
    .Y(_20576_));
 sky130_fd_sc_hd__nor2_1 _25421_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .Y(_20577_));
 sky130_vsdinv _25422_ (.A(\timer[19] ),
    .Y(_20578_));
 sky130_vsdinv _25423_ (.A(\timer[18] ),
    .Y(_20579_));
 sky130_fd_sc_hd__and3_1 _25424_ (.A(_20577_),
    .B(_20578_),
    .C(_20579_),
    .X(_20580_));
 sky130_fd_sc_hd__nand2_2 _25425_ (.A(_20576_),
    .B(_20580_),
    .Y(_20581_));
 sky130_fd_sc_hd__nor2_2 _25426_ (.A(_20556_),
    .B(_20581_),
    .Y(_20582_));
 sky130_fd_sc_hd__nor2_1 _25427_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .Y(_20583_));
 sky130_fd_sc_hd__nand2_1 _25428_ (.A(_20582_),
    .B(_20583_),
    .Y(_20584_));
 sky130_fd_sc_hd__or2_2 _25429_ (.A(\timer[26] ),
    .B(_20584_),
    .X(_20585_));
 sky130_fd_sc_hd__nor2_2 _25430_ (.A(\timer[27] ),
    .B(_20585_),
    .Y(_20586_));
 sky130_fd_sc_hd__nor2_1 _25431_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .Y(_20587_));
 sky130_fd_sc_hd__nand2_1 _25432_ (.A(_20586_),
    .B(_20587_),
    .Y(_20588_));
 sky130_fd_sc_hd__or2_4 _25433_ (.A(\timer[30] ),
    .B(_20588_),
    .X(_20589_));
 sky130_fd_sc_hd__nor2_8 _25434_ (.A(\timer[31] ),
    .B(_20589_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _25435_ (.A(\timer[0] ),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _25436_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .Y(_20590_));
 sky130_fd_sc_hd__nand2_1 _25437_ (.A(_20559_),
    .B(_20590_),
    .Y(_01211_));
 sky130_fd_sc_hd__and2_1 _25438_ (.A(_20559_),
    .B(\timer[2] ),
    .X(_20591_));
 sky130_fd_sc_hd__or2_1 _25439_ (.A(_20560_),
    .B(_20591_),
    .X(_01214_));
 sky130_fd_sc_hd__or2_1 _25440_ (.A(_20561_),
    .B(_20560_),
    .X(_20592_));
 sky130_fd_sc_hd__nand2_1 _25441_ (.A(_20592_),
    .B(_20562_),
    .Y(_01217_));
 sky130_fd_sc_hd__or2_1 _25442_ (.A(\timer[4] ),
    .B(_20562_),
    .X(_20593_));
 sky130_fd_sc_hd__nand2_1 _25443_ (.A(_20562_),
    .B(\timer[4] ),
    .Y(_20594_));
 sky130_fd_sc_hd__nand2_1 _25444_ (.A(_20593_),
    .B(_20594_),
    .Y(_01220_));
 sky130_fd_sc_hd__a21o_1 _25445_ (.A1(_20593_),
    .A2(\timer[5] ),
    .B1(_20563_),
    .X(_01223_));
 sky130_fd_sc_hd__nand2_1 _25446_ (.A(_20564_),
    .B(\timer[6] ),
    .Y(_20595_));
 sky130_fd_sc_hd__nand2_1 _25447_ (.A(_20566_),
    .B(_20595_),
    .Y(_01226_));
 sky130_vsdinv _25448_ (.A(\timer[7] ),
    .Y(_20596_));
 sky130_fd_sc_hd__nor2_1 _25449_ (.A(_20596_),
    .B(_20565_),
    .Y(_20597_));
 sky130_fd_sc_hd__or2_1 _25450_ (.A(_20597_),
    .B(_20567_),
    .X(_01229_));
 sky130_vsdinv _25451_ (.A(\timer[8] ),
    .Y(_20598_));
 sky130_fd_sc_hd__or2_1 _25452_ (.A(_20598_),
    .B(_20567_),
    .X(_20599_));
 sky130_fd_sc_hd__nand2_1 _25453_ (.A(_20567_),
    .B(_20598_),
    .Y(_20600_));
 sky130_fd_sc_hd__nand2_1 _25454_ (.A(_20599_),
    .B(_20600_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _25455_ (.A(_20600_),
    .B(\timer[9] ),
    .Y(_20601_));
 sky130_fd_sc_hd__nand2_1 _25456_ (.A(_20601_),
    .B(_20569_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand2_1 _25457_ (.A(_20569_),
    .B(\timer[10] ),
    .Y(_20602_));
 sky130_fd_sc_hd__nand2_1 _25458_ (.A(_20570_),
    .B(_20602_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _25459_ (.A(_20570_),
    .B(\timer[11] ),
    .Y(_20603_));
 sky130_fd_sc_hd__nand2_1 _25460_ (.A(_20571_),
    .B(_20603_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _25461_ (.A(_20571_),
    .B(\timer[12] ),
    .Y(_20604_));
 sky130_fd_sc_hd__nand2_1 _25462_ (.A(_20572_),
    .B(_20604_),
    .Y(_01244_));
 sky130_fd_sc_hd__and2_1 _25463_ (.A(_20572_),
    .B(\timer[13] ),
    .X(_20605_));
 sky130_fd_sc_hd__or2_1 _25464_ (.A(_20573_),
    .B(_20605_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_1 _25465_ (.A(_20574_),
    .B(_20573_),
    .X(_20606_));
 sky130_fd_sc_hd__nand2_1 _25466_ (.A(_20606_),
    .B(_20575_),
    .Y(_01250_));
 sky130_vsdinv _25467_ (.A(_20576_),
    .Y(_20607_));
 sky130_fd_sc_hd__nand2_1 _25468_ (.A(_20575_),
    .B(\timer[15] ),
    .Y(_20608_));
 sky130_fd_sc_hd__nand2_1 _25469_ (.A(_20607_),
    .B(_20608_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _25470_ (.A(_20607_),
    .B(\timer[16] ),
    .Y(_20609_));
 sky130_vsdinv _25471_ (.A(\timer[16] ),
    .Y(_20610_));
 sky130_fd_sc_hd__nand2_1 _25472_ (.A(_20576_),
    .B(_20610_),
    .Y(_20611_));
 sky130_fd_sc_hd__nand2_1 _25473_ (.A(_20609_),
    .B(_20611_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_1 _25474_ (.A(_20611_),
    .B(\timer[17] ),
    .Y(_20612_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(_20576_),
    .B(_20577_),
    .Y(_20613_));
 sky130_fd_sc_hd__nand2_1 _25476_ (.A(_20612_),
    .B(_20613_),
    .Y(_01259_));
 sky130_fd_sc_hd__or2_1 _25477_ (.A(\timer[18] ),
    .B(_20613_),
    .X(_20614_));
 sky130_fd_sc_hd__nand2_1 _25478_ (.A(_20613_),
    .B(\timer[18] ),
    .Y(_20615_));
 sky130_fd_sc_hd__nand2_1 _25479_ (.A(_20614_),
    .B(_20615_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_1 _25480_ (.A(_20614_),
    .B(\timer[19] ),
    .Y(_20616_));
 sky130_fd_sc_hd__nand2_1 _25481_ (.A(_20616_),
    .B(_20581_),
    .Y(_01265_));
 sky130_fd_sc_hd__or2_1 _25482_ (.A(\timer[20] ),
    .B(_20581_),
    .X(_20617_));
 sky130_fd_sc_hd__nand2_1 _25483_ (.A(_20581_),
    .B(\timer[20] ),
    .Y(_20618_));
 sky130_fd_sc_hd__nand2_1 _25484_ (.A(_20617_),
    .B(_20618_),
    .Y(_01268_));
 sky130_fd_sc_hd__or2_1 _25485_ (.A(\timer[21] ),
    .B(_20617_),
    .X(_20619_));
 sky130_fd_sc_hd__nand2_1 _25486_ (.A(_20617_),
    .B(\timer[21] ),
    .Y(_20620_));
 sky130_fd_sc_hd__nand2_1 _25487_ (.A(_20619_),
    .B(_20620_),
    .Y(_01271_));
 sky130_fd_sc_hd__or2_1 _25488_ (.A(\timer[22] ),
    .B(_20619_),
    .X(_20621_));
 sky130_fd_sc_hd__nand2_1 _25489_ (.A(_20619_),
    .B(\timer[22] ),
    .Y(_20622_));
 sky130_fd_sc_hd__nand2_1 _25490_ (.A(_20621_),
    .B(_20622_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2_1 _25491_ (.A(_20621_),
    .B(\timer[23] ),
    .Y(_20623_));
 sky130_vsdinv _25492_ (.A(_20582_),
    .Y(_20624_));
 sky130_fd_sc_hd__nand2_1 _25493_ (.A(_20623_),
    .B(_20624_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _25494_ (.A(_20624_),
    .B(\timer[24] ),
    .Y(_20625_));
 sky130_vsdinv _25495_ (.A(\timer[24] ),
    .Y(_20626_));
 sky130_fd_sc_hd__nand2_1 _25496_ (.A(_20582_),
    .B(_20626_),
    .Y(_20627_));
 sky130_fd_sc_hd__nand2_1 _25497_ (.A(_20625_),
    .B(_20627_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_1 _25498_ (.A(_20627_),
    .B(\timer[25] ),
    .Y(_20628_));
 sky130_fd_sc_hd__nand2_1 _25499_ (.A(_20628_),
    .B(_20584_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_1 _25500_ (.A(_20584_),
    .B(\timer[26] ),
    .Y(_20629_));
 sky130_fd_sc_hd__nand2_1 _25501_ (.A(_20585_),
    .B(_20629_),
    .Y(_01286_));
 sky130_vsdinv _25502_ (.A(_20586_),
    .Y(_20630_));
 sky130_fd_sc_hd__nand2_1 _25503_ (.A(_20585_),
    .B(\timer[27] ),
    .Y(_20631_));
 sky130_fd_sc_hd__nand2_1 _25504_ (.A(_20630_),
    .B(_20631_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_1 _25505_ (.A(_20630_),
    .B(\timer[28] ),
    .Y(_20632_));
 sky130_vsdinv _25506_ (.A(\timer[28] ),
    .Y(_20633_));
 sky130_fd_sc_hd__nand2_1 _25507_ (.A(_20586_),
    .B(_20633_),
    .Y(_20634_));
 sky130_fd_sc_hd__nand2_1 _25508_ (.A(_20632_),
    .B(_20634_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _25509_ (.A(_20634_),
    .B(\timer[29] ),
    .Y(_20635_));
 sky130_fd_sc_hd__nand2_1 _25510_ (.A(_20635_),
    .B(_20588_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _25511_ (.A(_20588_),
    .B(\timer[30] ),
    .Y(_20636_));
 sky130_fd_sc_hd__nand2_1 _25512_ (.A(_20589_),
    .B(_20636_),
    .Y(_01298_));
 sky130_fd_sc_hd__and2_1 _25513_ (.A(_20589_),
    .B(\timer[31] ),
    .X(_20637_));
 sky130_fd_sc_hd__or2_1 _25514_ (.A(_01208_),
    .B(_20637_),
    .X(_01301_));
 sky130_fd_sc_hd__clkbuf_2 _25515_ (.A(_19958_),
    .X(_20638_));
 sky130_vsdinv _25516_ (.A(\decoded_imm[5] ),
    .Y(_20639_));
 sky130_fd_sc_hd__nor2_1 _25517_ (.A(_20638_),
    .B(_20639_),
    .Y(_01315_));
 sky130_vsdinv _25518_ (.A(\decoded_imm[6] ),
    .Y(_20640_));
 sky130_fd_sc_hd__nor2_1 _25519_ (.A(_20638_),
    .B(_20640_),
    .Y(_01317_));
 sky130_vsdinv _25520_ (.A(\decoded_imm[7] ),
    .Y(_20641_));
 sky130_fd_sc_hd__nor2_1 _25521_ (.A(_20638_),
    .B(_20641_),
    .Y(_01319_));
 sky130_vsdinv _25522_ (.A(\decoded_imm[8] ),
    .Y(_20642_));
 sky130_fd_sc_hd__nor2_1 _25523_ (.A(_20638_),
    .B(_20642_),
    .Y(_01321_));
 sky130_vsdinv _25524_ (.A(\decoded_imm[9] ),
    .Y(_20643_));
 sky130_fd_sc_hd__nor2_1 _25525_ (.A(_20638_),
    .B(_20643_),
    .Y(_01323_));
 sky130_fd_sc_hd__clkbuf_2 _25526_ (.A(_19958_),
    .X(_20644_));
 sky130_vsdinv _25527_ (.A(\decoded_imm[10] ),
    .Y(_20645_));
 sky130_fd_sc_hd__nor2_1 _25528_ (.A(_20644_),
    .B(_20645_),
    .Y(_01325_));
 sky130_vsdinv _25529_ (.A(\decoded_imm[11] ),
    .Y(_20646_));
 sky130_fd_sc_hd__nor2_1 _25530_ (.A(_20644_),
    .B(_20646_),
    .Y(_01327_));
 sky130_vsdinv _25531_ (.A(\decoded_imm[12] ),
    .Y(_20647_));
 sky130_fd_sc_hd__nor2_1 _25532_ (.A(_20644_),
    .B(_20647_),
    .Y(_01329_));
 sky130_vsdinv _25533_ (.A(\decoded_imm[13] ),
    .Y(_20648_));
 sky130_fd_sc_hd__nor2_1 _25534_ (.A(_20644_),
    .B(_20648_),
    .Y(_01331_));
 sky130_vsdinv _25535_ (.A(\decoded_imm[14] ),
    .Y(_20649_));
 sky130_fd_sc_hd__nor2_1 _25536_ (.A(_20644_),
    .B(_20649_),
    .Y(_01333_));
 sky130_vsdinv _25537_ (.A(\decoded_imm[15] ),
    .Y(_20650_));
 sky130_fd_sc_hd__nor2_1 _25538_ (.A(_20644_),
    .B(_20650_),
    .Y(_01335_));
 sky130_fd_sc_hd__clkbuf_2 _25539_ (.A(is_slli_srli_srai),
    .X(_20651_));
 sky130_vsdinv _25540_ (.A(\decoded_imm[16] ),
    .Y(_20652_));
 sky130_fd_sc_hd__nor2_1 _25541_ (.A(_20651_),
    .B(_20652_),
    .Y(_01337_));
 sky130_vsdinv _25542_ (.A(\decoded_imm[17] ),
    .Y(_20653_));
 sky130_fd_sc_hd__nor2_1 _25543_ (.A(_20651_),
    .B(_20653_),
    .Y(_01339_));
 sky130_vsdinv _25544_ (.A(\decoded_imm[18] ),
    .Y(_20654_));
 sky130_fd_sc_hd__nor2_1 _25545_ (.A(_20651_),
    .B(_20654_),
    .Y(_01341_));
 sky130_vsdinv _25546_ (.A(\decoded_imm[19] ),
    .Y(_20655_));
 sky130_fd_sc_hd__nor2_1 _25547_ (.A(_20651_),
    .B(_20655_),
    .Y(_01343_));
 sky130_vsdinv _25548_ (.A(\decoded_imm[20] ),
    .Y(_20656_));
 sky130_fd_sc_hd__nor2_1 _25549_ (.A(_20651_),
    .B(_20656_),
    .Y(_01345_));
 sky130_fd_sc_hd__inv_2 _25550_ (.A(\decoded_imm[21] ),
    .Y(_20657_));
 sky130_fd_sc_hd__nor2_1 _25551_ (.A(_20651_),
    .B(_20657_),
    .Y(_01347_));
 sky130_fd_sc_hd__buf_2 _25552_ (.A(is_slli_srli_srai),
    .X(_20658_));
 sky130_vsdinv _25553_ (.A(\decoded_imm[22] ),
    .Y(_20659_));
 sky130_fd_sc_hd__nor2_1 _25554_ (.A(_20658_),
    .B(_20659_),
    .Y(_01349_));
 sky130_vsdinv _25555_ (.A(\decoded_imm[23] ),
    .Y(_20660_));
 sky130_fd_sc_hd__nor2_1 _25556_ (.A(_20658_),
    .B(_20660_),
    .Y(_01351_));
 sky130_vsdinv _25557_ (.A(\decoded_imm[24] ),
    .Y(_20661_));
 sky130_fd_sc_hd__nor2_1 _25558_ (.A(_20658_),
    .B(_20661_),
    .Y(_01353_));
 sky130_vsdinv _25559_ (.A(\decoded_imm[25] ),
    .Y(_20662_));
 sky130_fd_sc_hd__nor2_1 _25560_ (.A(_20658_),
    .B(_20662_),
    .Y(_01355_));
 sky130_fd_sc_hd__inv_2 _25561_ (.A(\decoded_imm[26] ),
    .Y(_20663_));
 sky130_fd_sc_hd__nor2_1 _25562_ (.A(_20658_),
    .B(_20663_),
    .Y(_01357_));
 sky130_vsdinv _25563_ (.A(\decoded_imm[27] ),
    .Y(_20664_));
 sky130_fd_sc_hd__nor2_1 _25564_ (.A(_20658_),
    .B(_20664_),
    .Y(_01359_));
 sky130_vsdinv _25565_ (.A(\decoded_imm[28] ),
    .Y(_20665_));
 sky130_fd_sc_hd__nor2_1 _25566_ (.A(_19958_),
    .B(_20665_),
    .Y(_01361_));
 sky130_fd_sc_hd__inv_2 _25567_ (.A(\decoded_imm[29] ),
    .Y(_20666_));
 sky130_fd_sc_hd__nor2_1 _25568_ (.A(_19958_),
    .B(_20666_),
    .Y(_01363_));
 sky130_vsdinv _25569_ (.A(\decoded_imm[30] ),
    .Y(_20667_));
 sky130_fd_sc_hd__nor2_1 _25570_ (.A(_19958_),
    .B(_20667_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2b_1 _25571_ (.A(_20638_),
    .B_N(\decoded_imm[31] ),
    .Y(_01367_));
 sky130_fd_sc_hd__clkbuf_2 _25572_ (.A(_20023_),
    .X(_20668_));
 sky130_vsdinv _25573_ (.A(\reg_next_pc[0] ),
    .Y(_20669_));
 sky130_fd_sc_hd__nor2_1 _25574_ (.A(_20668_),
    .B(_20669_),
    .Y(_01369_));
 sky130_vsdinv _25575_ (.A(\decoded_imm[0] ),
    .Y(_20670_));
 sky130_fd_sc_hd__nand2_1 _25576_ (.A(_20670_),
    .B(_20323_),
    .Y(_20671_));
 sky130_fd_sc_hd__nand2_1 _25577_ (.A(\decoded_imm[0] ),
    .B(net306),
    .Y(_20672_));
 sky130_fd_sc_hd__and2_1 _25578_ (.A(_20671_),
    .B(_20672_),
    .X(_01371_));
 sky130_fd_sc_hd__nor2_1 _25579_ (.A(_20668_),
    .B(_19091_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _25580_ (.A(net317),
    .B(\decoded_imm[1] ),
    .Y(_20673_));
 sky130_fd_sc_hd__nand2_1 _25581_ (.A(net317),
    .B(\decoded_imm[1] ),
    .Y(_20674_));
 sky130_fd_sc_hd__or2b_1 _25582_ (.A(_20673_),
    .B_N(_20674_),
    .X(_20675_));
 sky130_fd_sc_hd__xor2_1 _25583_ (.A(_20672_),
    .B(_20675_),
    .X(_01374_));
 sky130_fd_sc_hd__inv_2 _25584_ (.A(\reg_pc[2] ),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _25585_ (.A(_20668_),
    .B(_02073_),
    .Y(_01375_));
 sky130_fd_sc_hd__o21ai_1 _25586_ (.A1(_20672_),
    .A2(_20673_),
    .B1(_20674_),
    .Y(_20676_));
 sky130_fd_sc_hd__xnor2_1 _25587_ (.A(_20062_),
    .B(\decoded_imm[2] ),
    .Y(_20677_));
 sky130_fd_sc_hd__xnor2_1 _25588_ (.A(_20676_),
    .B(_20677_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _25589_ (.A(_20668_),
    .B(_19087_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _25590_ (.A(net331),
    .B(\decoded_imm[3] ),
    .Y(_20678_));
 sky130_fd_sc_hd__nand2_1 _25591_ (.A(net331),
    .B(\decoded_imm[3] ),
    .Y(_20679_));
 sky130_fd_sc_hd__or2b_1 _25592_ (.A(_20678_),
    .B_N(_20679_),
    .X(_20680_));
 sky130_fd_sc_hd__o21ai_1 _25593_ (.A1(_20062_),
    .A2(\decoded_imm[2] ),
    .B1(_20676_),
    .Y(_20681_));
 sky130_fd_sc_hd__o21a_1 _25594_ (.A1(_20482_),
    .A2(_20240_),
    .B1(_20681_),
    .X(_20682_));
 sky130_fd_sc_hd__xor2_1 _25595_ (.A(_20680_),
    .B(_20682_),
    .X(_01380_));
 sky130_vsdinv _25596_ (.A(\reg_pc[4] ),
    .Y(_20683_));
 sky130_fd_sc_hd__nor2_1 _25597_ (.A(_20668_),
    .B(_20683_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _25598_ (.A(net332),
    .B(\decoded_imm[4] ),
    .Y(_20684_));
 sky130_fd_sc_hd__nor2_1 _25599_ (.A(_20488_),
    .B(_20250_),
    .Y(_20685_));
 sky130_fd_sc_hd__nor2_1 _25600_ (.A(_20684_),
    .B(_20685_),
    .Y(_20686_));
 sky130_fd_sc_hd__o21ai_2 _25601_ (.A1(_20678_),
    .A2(_20682_),
    .B1(_20679_),
    .Y(_20687_));
 sky130_fd_sc_hd__xor2_1 _25602_ (.A(_20686_),
    .B(_20687_),
    .X(_01383_));
 sky130_vsdinv _25603_ (.A(\reg_pc[5] ),
    .Y(_20688_));
 sky130_fd_sc_hd__nor2_1 _25604_ (.A(_20668_),
    .B(_20688_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _25605_ (.A(_20059_),
    .B(\decoded_imm[5] ),
    .Y(_20689_));
 sky130_fd_sc_hd__nor2_2 _25606_ (.A(_20469_),
    .B(_20639_),
    .Y(_20690_));
 sky130_fd_sc_hd__or2_1 _25607_ (.A(_20689_),
    .B(_20690_),
    .X(_20691_));
 sky130_vsdinv _25608_ (.A(_20684_),
    .Y(_20692_));
 sky130_fd_sc_hd__a21oi_2 _25609_ (.A1(_20687_),
    .A2(_20692_),
    .B1(_20685_),
    .Y(_20693_));
 sky130_fd_sc_hd__xor2_1 _25610_ (.A(_20691_),
    .B(_20693_),
    .X(_01386_));
 sky130_fd_sc_hd__clkbuf_2 _25611_ (.A(_20023_),
    .X(_20694_));
 sky130_vsdinv _25612_ (.A(\reg_pc[6] ),
    .Y(_20695_));
 sky130_fd_sc_hd__nor2_1 _25613_ (.A(_20694_),
    .B(_20695_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_1 _25614_ (.A(net334),
    .B(\decoded_imm[6] ),
    .X(_20696_));
 sky130_fd_sc_hd__nor2_1 _25615_ (.A(_20689_),
    .B(_20693_),
    .Y(_20697_));
 sky130_fd_sc_hd__or2_1 _25616_ (.A(_20690_),
    .B(_20697_),
    .X(_20698_));
 sky130_fd_sc_hd__or2_1 _25617_ (.A(_20696_),
    .B(_20698_),
    .X(_20699_));
 sky130_fd_sc_hd__nand2_1 _25618_ (.A(_20698_),
    .B(_20696_),
    .Y(_20700_));
 sky130_fd_sc_hd__and2_1 _25619_ (.A(_20699_),
    .B(_20700_),
    .X(_01389_));
 sky130_vsdinv _25620_ (.A(\reg_pc[7] ),
    .Y(_20701_));
 sky130_fd_sc_hd__nor2_1 _25621_ (.A(_20694_),
    .B(_20701_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_1 _25622_ (.A(_20057_),
    .B(\decoded_imm[7] ),
    .Y(_20702_));
 sky130_vsdinv _25623_ (.A(net335),
    .Y(_20703_));
 sky130_fd_sc_hd__nor2_1 _25624_ (.A(_20703_),
    .B(_20641_),
    .Y(_20704_));
 sky130_fd_sc_hd__nor2_1 _25625_ (.A(_20702_),
    .B(_20704_),
    .Y(_20705_));
 sky130_fd_sc_hd__o21ai_1 _25626_ (.A1(_20472_),
    .A2(_20640_),
    .B1(_20700_),
    .Y(_20706_));
 sky130_fd_sc_hd__xor2_1 _25627_ (.A(_20705_),
    .B(_20706_),
    .X(_01392_));
 sky130_vsdinv _25628_ (.A(\reg_pc[8] ),
    .Y(_20707_));
 sky130_fd_sc_hd__nor2_1 _25629_ (.A(_20694_),
    .B(_20707_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _25630_ (.A(net336),
    .B(\decoded_imm[8] ),
    .Y(_20708_));
 sky130_fd_sc_hd__nor2_1 _25631_ (.A(_20460_),
    .B(_20642_),
    .Y(_20709_));
 sky130_fd_sc_hd__nor2_1 _25632_ (.A(_20708_),
    .B(_20709_),
    .Y(_20710_));
 sky130_fd_sc_hd__and2_1 _25633_ (.A(_20705_),
    .B(_20696_),
    .X(_20711_));
 sky130_fd_sc_hd__o21ai_2 _25634_ (.A1(_20690_),
    .A2(_20697_),
    .B1(_20711_),
    .Y(_20712_));
 sky130_vsdinv _25635_ (.A(_20704_),
    .Y(_20713_));
 sky130_fd_sc_hd__o31a_1 _25636_ (.A1(_20472_),
    .A2(_20640_),
    .A3(_20702_),
    .B1(_20713_),
    .X(_20714_));
 sky130_fd_sc_hd__nand2_1 _25637_ (.A(_20712_),
    .B(_20714_),
    .Y(_20715_));
 sky130_fd_sc_hd__xor2_1 _25638_ (.A(_20710_),
    .B(_20715_),
    .X(_01395_));
 sky130_vsdinv _25639_ (.A(\reg_pc[9] ),
    .Y(_20716_));
 sky130_fd_sc_hd__nor2_1 _25640_ (.A(_20694_),
    .B(_20716_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _25641_ (.A(_20055_),
    .B(\decoded_imm[9] ),
    .Y(_20717_));
 sky130_fd_sc_hd__nor2_1 _25642_ (.A(_20456_),
    .B(_20643_),
    .Y(_20718_));
 sky130_fd_sc_hd__nor2_2 _25643_ (.A(_20717_),
    .B(_20718_),
    .Y(_20719_));
 sky130_vsdinv _25644_ (.A(_20715_),
    .Y(_20720_));
 sky130_fd_sc_hd__o21ba_1 _25645_ (.A1(_20708_),
    .A2(_20720_),
    .B1_N(_20709_),
    .X(_20721_));
 sky130_fd_sc_hd__xnor2_1 _25646_ (.A(_20719_),
    .B(_20721_),
    .Y(_01398_));
 sky130_vsdinv _25647_ (.A(\reg_pc[10] ),
    .Y(_20722_));
 sky130_fd_sc_hd__nor2_1 _25648_ (.A(_20694_),
    .B(_20722_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_1 _25649_ (.A(_20054_),
    .B(\decoded_imm[10] ),
    .Y(_20723_));
 sky130_fd_sc_hd__nor2_1 _25650_ (.A(_20464_),
    .B(_20645_),
    .Y(_20724_));
 sky130_fd_sc_hd__nor2_1 _25651_ (.A(_20723_),
    .B(_20724_),
    .Y(_20725_));
 sky130_vsdinv _25652_ (.A(_20717_),
    .Y(_20726_));
 sky130_fd_sc_hd__a21o_1 _25653_ (.A1(_20709_),
    .A2(_20726_),
    .B1(_20718_),
    .X(_20727_));
 sky130_fd_sc_hd__nand2_1 _25654_ (.A(_20710_),
    .B(_20719_),
    .Y(_20728_));
 sky130_fd_sc_hd__a21oi_2 _25655_ (.A1(_20712_),
    .A2(_20714_),
    .B1(_20728_),
    .Y(_20729_));
 sky130_fd_sc_hd__nor3_1 _25656_ (.A(_20725_),
    .B(_20727_),
    .C(_20729_),
    .Y(_20730_));
 sky130_fd_sc_hd__o21ai_2 _25657_ (.A1(_20727_),
    .A2(_20729_),
    .B1(_20725_),
    .Y(_20731_));
 sky130_fd_sc_hd__nor2b_1 _25658_ (.A(_20730_),
    .B_N(_20731_),
    .Y(_01401_));
 sky130_vsdinv _25659_ (.A(\reg_pc[11] ),
    .Y(_20732_));
 sky130_fd_sc_hd__nor2_1 _25660_ (.A(_20694_),
    .B(_20732_),
    .Y(_01402_));
 sky130_vsdinv _25661_ (.A(_20724_),
    .Y(_20733_));
 sky130_fd_sc_hd__nor2_1 _25662_ (.A(net308),
    .B(\decoded_imm[11] ),
    .Y(_20734_));
 sky130_fd_sc_hd__nor2_2 _25663_ (.A(_20452_),
    .B(_20646_),
    .Y(_20735_));
 sky130_fd_sc_hd__or2_1 _25664_ (.A(_20734_),
    .B(_20735_),
    .X(_20736_));
 sky130_fd_sc_hd__a21oi_2 _25665_ (.A1(_20731_),
    .A2(_20733_),
    .B1(_20736_),
    .Y(_20737_));
 sky130_fd_sc_hd__and3_1 _25666_ (.A(_20731_),
    .B(_20733_),
    .C(_20736_),
    .X(_20738_));
 sky130_fd_sc_hd__nor2_1 _25667_ (.A(_20737_),
    .B(_20738_),
    .Y(_01404_));
 sky130_fd_sc_hd__buf_2 _25668_ (.A(_20023_),
    .X(_20739_));
 sky130_vsdinv _25669_ (.A(\reg_pc[12] ),
    .Y(_20740_));
 sky130_fd_sc_hd__nor2_1 _25670_ (.A(_20739_),
    .B(_20740_),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _25671_ (.A(net309),
    .B(_20647_),
    .Y(_20741_));
 sky130_fd_sc_hd__nor2_1 _25672_ (.A(\decoded_imm[12] ),
    .B(_20436_),
    .Y(_20742_));
 sky130_fd_sc_hd__or4_1 _25673_ (.A(_20735_),
    .B(_20741_),
    .C(_20742_),
    .D(_20737_),
    .X(_20743_));
 sky130_fd_sc_hd__nor2_1 _25674_ (.A(_20741_),
    .B(_20742_),
    .Y(_20744_));
 sky130_fd_sc_hd__o21bai_2 _25675_ (.A1(_20735_),
    .A2(_20737_),
    .B1_N(_20744_),
    .Y(_20745_));
 sky130_fd_sc_hd__and2_1 _25676_ (.A(_20743_),
    .B(_20745_),
    .X(_01407_));
 sky130_vsdinv _25677_ (.A(\reg_pc[13] ),
    .Y(_20746_));
 sky130_fd_sc_hd__nor2_1 _25678_ (.A(_20739_),
    .B(_20746_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_1 _25679_ (.A(_20436_),
    .B(_20647_),
    .Y(_20747_));
 sky130_vsdinv _25680_ (.A(_20747_),
    .Y(_20748_));
 sky130_fd_sc_hd__nor2_1 _25681_ (.A(net310),
    .B(\decoded_imm[13] ),
    .Y(_20749_));
 sky130_fd_sc_hd__nor2_2 _25682_ (.A(_20431_),
    .B(_20648_),
    .Y(_20750_));
 sky130_fd_sc_hd__or2_2 _25683_ (.A(_20749_),
    .B(_20750_),
    .X(_20751_));
 sky130_fd_sc_hd__a21oi_4 _25684_ (.A1(_20745_),
    .A2(_20748_),
    .B1(_20751_),
    .Y(_20752_));
 sky130_fd_sc_hd__and3_1 _25685_ (.A(_20745_),
    .B(_20748_),
    .C(_20751_),
    .X(_20753_));
 sky130_fd_sc_hd__nor2_1 _25686_ (.A(_20752_),
    .B(_20753_),
    .Y(_01410_));
 sky130_vsdinv _25687_ (.A(\reg_pc[14] ),
    .Y(_20754_));
 sky130_fd_sc_hd__nor2_1 _25688_ (.A(_20739_),
    .B(_20754_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_2 _25689_ (.A(net311),
    .B(_20649_),
    .Y(_20755_));
 sky130_fd_sc_hd__nor2_2 _25690_ (.A(\decoded_imm[14] ),
    .B(_20441_),
    .Y(_20756_));
 sky130_fd_sc_hd__or4_1 _25691_ (.A(_20750_),
    .B(_20755_),
    .C(_20756_),
    .D(_20752_),
    .X(_20757_));
 sky130_fd_sc_hd__o22ai_4 _25692_ (.A1(_20755_),
    .A2(_20756_),
    .B1(_20750_),
    .B2(_20752_),
    .Y(_20758_));
 sky130_fd_sc_hd__and2_1 _25693_ (.A(_20757_),
    .B(_20758_),
    .X(_01413_));
 sky130_vsdinv _25694_ (.A(\reg_pc[15] ),
    .Y(_20759_));
 sky130_fd_sc_hd__nor2_1 _25695_ (.A(_20739_),
    .B(_20759_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _25696_ (.A(_20441_),
    .B(_20649_),
    .Y(_20760_));
 sky130_vsdinv _25697_ (.A(_20760_),
    .Y(_20761_));
 sky130_fd_sc_hd__nor2_1 _25698_ (.A(net312),
    .B(\decoded_imm[15] ),
    .Y(_20762_));
 sky130_fd_sc_hd__nor2_4 _25699_ (.A(_20445_),
    .B(_20650_),
    .Y(_20763_));
 sky130_fd_sc_hd__nor2_1 _25700_ (.A(_20762_),
    .B(_20763_),
    .Y(_20764_));
 sky130_fd_sc_hd__a21boi_4 _25701_ (.A1(_20758_),
    .A2(_20761_),
    .B1_N(_20764_),
    .Y(_20765_));
 sky130_fd_sc_hd__o211a_1 _25702_ (.A1(_20763_),
    .A2(_20762_),
    .B1(_20761_),
    .C1(_20758_),
    .X(_20766_));
 sky130_fd_sc_hd__nor2_1 _25703_ (.A(_20765_),
    .B(_20766_),
    .Y(_01416_));
 sky130_vsdinv _25704_ (.A(\reg_pc[16] ),
    .Y(_20767_));
 sky130_fd_sc_hd__nor2_1 _25705_ (.A(_20739_),
    .B(_20767_),
    .Y(_01417_));
 sky130_fd_sc_hd__xnor2_1 _25706_ (.A(_20050_),
    .B(\decoded_imm[16] ),
    .Y(_20768_));
 sky130_fd_sc_hd__nor2_1 _25707_ (.A(_20763_),
    .B(_20765_),
    .Y(_20769_));
 sky130_fd_sc_hd__or2_1 _25708_ (.A(_20768_),
    .B(_20769_),
    .X(_20770_));
 sky130_fd_sc_hd__nand2_1 _25709_ (.A(_20769_),
    .B(_20768_),
    .Y(_20771_));
 sky130_fd_sc_hd__and2_1 _25710_ (.A(_20770_),
    .B(_20771_),
    .X(_01419_));
 sky130_vsdinv _25711_ (.A(\reg_pc[17] ),
    .Y(_20772_));
 sky130_fd_sc_hd__nor2_1 _25712_ (.A(_20739_),
    .B(_20772_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _25713_ (.A(net314),
    .B(\decoded_imm[17] ),
    .Y(_20773_));
 sky130_fd_sc_hd__nor2_1 _25714_ (.A(_20396_),
    .B(_20653_),
    .Y(_20774_));
 sky130_fd_sc_hd__nor2_1 _25715_ (.A(_20773_),
    .B(_20774_),
    .Y(_20775_));
 sky130_fd_sc_hd__inv_2 _25716_ (.A(net313),
    .Y(_20776_));
 sky130_fd_sc_hd__o21ai_1 _25717_ (.A1(_20776_),
    .A2(_20652_),
    .B1(_20770_),
    .Y(_20777_));
 sky130_fd_sc_hd__xor2_1 _25718_ (.A(_20775_),
    .B(_20777_),
    .X(_01422_));
 sky130_fd_sc_hd__buf_2 _25719_ (.A(instr_lui),
    .X(_20778_));
 sky130_vsdinv _25720_ (.A(\reg_pc[18] ),
    .Y(_20779_));
 sky130_fd_sc_hd__nor2_1 _25721_ (.A(_20778_),
    .B(_20779_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _25722_ (.A(_20049_),
    .B(\decoded_imm[18] ),
    .Y(_20780_));
 sky130_fd_sc_hd__nor2_4 _25723_ (.A(_20404_),
    .B(_20654_),
    .Y(_20781_));
 sky130_fd_sc_hd__nor2_1 _25724_ (.A(_20780_),
    .B(_20781_),
    .Y(_20782_));
 sky130_fd_sc_hd__and2b_1 _25725_ (.A_N(_20768_),
    .B(_20775_),
    .X(_20783_));
 sky130_fd_sc_hd__o21ai_2 _25726_ (.A1(_20763_),
    .A2(_20765_),
    .B1(_20783_),
    .Y(_20784_));
 sky130_vsdinv _25727_ (.A(_20774_),
    .Y(_20785_));
 sky130_fd_sc_hd__o31a_1 _25728_ (.A1(_20776_),
    .A2(_20652_),
    .A3(_20773_),
    .B1(_20785_),
    .X(_20786_));
 sky130_fd_sc_hd__nand2_1 _25729_ (.A(_20784_),
    .B(_20786_),
    .Y(_20787_));
 sky130_fd_sc_hd__xor2_1 _25730_ (.A(_20782_),
    .B(_20787_),
    .X(_01425_));
 sky130_vsdinv _25731_ (.A(\reg_pc[19] ),
    .Y(_20788_));
 sky130_fd_sc_hd__nor2_1 _25732_ (.A(_20778_),
    .B(_20788_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_2 _25733_ (.A(_20047_),
    .B(_20655_),
    .Y(_20789_));
 sky130_fd_sc_hd__nor2_2 _25734_ (.A(\decoded_imm[19] ),
    .B(_20400_),
    .Y(_20790_));
 sky130_fd_sc_hd__a22oi_4 _25735_ (.A1(_20404_),
    .A2(_20654_),
    .B1(_20784_),
    .B2(_20786_),
    .Y(_20791_));
 sky130_fd_sc_hd__or4_1 _25736_ (.A(_20781_),
    .B(_20789_),
    .C(_20790_),
    .D(_20791_),
    .X(_20792_));
 sky130_fd_sc_hd__o22ai_4 _25737_ (.A1(_20789_),
    .A2(_20790_),
    .B1(_20781_),
    .B2(_20791_),
    .Y(_20793_));
 sky130_fd_sc_hd__and2_1 _25738_ (.A(_20792_),
    .B(_20793_),
    .X(_01428_));
 sky130_vsdinv _25739_ (.A(\reg_pc[20] ),
    .Y(_20794_));
 sky130_fd_sc_hd__nor2_1 _25740_ (.A(_20778_),
    .B(_20794_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_2 _25741_ (.A(_20047_),
    .B(\decoded_imm[19] ),
    .Y(_20795_));
 sky130_fd_sc_hd__nor2_1 _25742_ (.A(_20046_),
    .B(\decoded_imm[20] ),
    .Y(_20796_));
 sky130_fd_sc_hd__nor2_4 _25743_ (.A(_20423_),
    .B(_20656_),
    .Y(_20797_));
 sky130_fd_sc_hd__nor2_1 _25744_ (.A(_20796_),
    .B(_20797_),
    .Y(_20798_));
 sky130_vsdinv _25745_ (.A(_20798_),
    .Y(_20799_));
 sky130_fd_sc_hd__a21oi_4 _25746_ (.A1(_20793_),
    .A2(_20795_),
    .B1(_20799_),
    .Y(_20800_));
 sky130_fd_sc_hd__and3_1 _25747_ (.A(_20793_),
    .B(_20795_),
    .C(_20799_),
    .X(_20801_));
 sky130_fd_sc_hd__nor2_1 _25748_ (.A(_20800_),
    .B(_20801_),
    .Y(_01431_));
 sky130_vsdinv _25749_ (.A(\reg_pc[21] ),
    .Y(_20802_));
 sky130_fd_sc_hd__nor2_1 _25750_ (.A(_20778_),
    .B(_20802_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_2 _25751_ (.A(_20045_),
    .B(_20657_),
    .Y(_20803_));
 sky130_fd_sc_hd__nor2_2 _25752_ (.A(\decoded_imm[21] ),
    .B(_20415_),
    .Y(_20804_));
 sky130_fd_sc_hd__or4_1 _25753_ (.A(_20797_),
    .B(_20803_),
    .C(_20804_),
    .D(_20800_),
    .X(_20805_));
 sky130_fd_sc_hd__o22ai_4 _25754_ (.A1(_20803_),
    .A2(_20804_),
    .B1(_20797_),
    .B2(_20800_),
    .Y(_20806_));
 sky130_fd_sc_hd__and2_1 _25755_ (.A(_20805_),
    .B(_20806_),
    .X(_01434_));
 sky130_vsdinv _25756_ (.A(\reg_pc[22] ),
    .Y(_20807_));
 sky130_fd_sc_hd__nor2_1 _25757_ (.A(_20778_),
    .B(_20807_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_2 _25758_ (.A(_20045_),
    .B(\decoded_imm[21] ),
    .Y(_20808_));
 sky130_fd_sc_hd__nor2_1 _25759_ (.A(_20044_),
    .B(\decoded_imm[22] ),
    .Y(_20809_));
 sky130_fd_sc_hd__nor2_4 _25760_ (.A(_20411_),
    .B(_20659_),
    .Y(_20810_));
 sky130_fd_sc_hd__nor2_1 _25761_ (.A(_20809_),
    .B(_20810_),
    .Y(_20811_));
 sky130_vsdinv _25762_ (.A(_20811_),
    .Y(_20812_));
 sky130_fd_sc_hd__a21oi_4 _25763_ (.A1(_20806_),
    .A2(_20808_),
    .B1(_20812_),
    .Y(_20813_));
 sky130_fd_sc_hd__and3_1 _25764_ (.A(_20806_),
    .B(_20808_),
    .C(_20812_),
    .X(_20814_));
 sky130_fd_sc_hd__nor2_1 _25765_ (.A(_20813_),
    .B(_20814_),
    .Y(_01437_));
 sky130_vsdinv _25766_ (.A(\reg_pc[23] ),
    .Y(_20815_));
 sky130_fd_sc_hd__nor2_2 _25767_ (.A(_20778_),
    .B(_20815_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_2 _25768_ (.A(_20043_),
    .B(_20660_),
    .Y(_20816_));
 sky130_fd_sc_hd__nor2_2 _25769_ (.A(\decoded_imm[23] ),
    .B(_20418_),
    .Y(_20817_));
 sky130_fd_sc_hd__or4_1 _25770_ (.A(_20810_),
    .B(_20816_),
    .C(_20817_),
    .D(_20813_),
    .X(_20818_));
 sky130_fd_sc_hd__o22ai_4 _25771_ (.A1(_20816_),
    .A2(_20817_),
    .B1(_20810_),
    .B2(_20813_),
    .Y(_20819_));
 sky130_fd_sc_hd__and2_1 _25772_ (.A(_20818_),
    .B(_20819_),
    .X(_01440_));
 sky130_fd_sc_hd__clkbuf_2 _25773_ (.A(instr_lui),
    .X(_20820_));
 sky130_vsdinv _25774_ (.A(\reg_pc[24] ),
    .Y(_20821_));
 sky130_fd_sc_hd__nor2_2 _25775_ (.A(_20820_),
    .B(_20821_),
    .Y(_01441_));
 sky130_fd_sc_hd__xor2_2 _25776_ (.A(_20042_),
    .B(\decoded_imm[24] ),
    .X(_20822_));
 sky130_fd_sc_hd__nand2_2 _25777_ (.A(_20043_),
    .B(\decoded_imm[23] ),
    .Y(_20823_));
 sky130_fd_sc_hd__nand2_1 _25778_ (.A(_20819_),
    .B(_20823_),
    .Y(_20824_));
 sky130_fd_sc_hd__or2_1 _25779_ (.A(_20822_),
    .B(_20824_),
    .X(_20825_));
 sky130_fd_sc_hd__nand2_1 _25780_ (.A(_20824_),
    .B(_20822_),
    .Y(_20826_));
 sky130_fd_sc_hd__and2_1 _25781_ (.A(_20825_),
    .B(_20826_),
    .X(_01443_));
 sky130_vsdinv _25782_ (.A(\reg_pc[25] ),
    .Y(_20827_));
 sky130_fd_sc_hd__nor2_1 _25783_ (.A(_20820_),
    .B(_20827_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _25784_ (.A(_20040_),
    .B(\decoded_imm[25] ),
    .Y(_20828_));
 sky130_fd_sc_hd__nor2_1 _25785_ (.A(_20501_),
    .B(_20662_),
    .Y(_20829_));
 sky130_fd_sc_hd__or2_1 _25786_ (.A(_20828_),
    .B(_20829_),
    .X(_20830_));
 sky130_vsdinv _25787_ (.A(_20830_),
    .Y(_20831_));
 sky130_fd_sc_hd__o21ai_1 _25788_ (.A1(_20513_),
    .A2(_20661_),
    .B1(_20826_),
    .Y(_20832_));
 sky130_fd_sc_hd__xor2_1 _25789_ (.A(_20831_),
    .B(_20832_),
    .X(_01446_));
 sky130_vsdinv _25790_ (.A(\reg_pc[26] ),
    .Y(_20833_));
 sky130_fd_sc_hd__nor2_1 _25791_ (.A(_20820_),
    .B(_20833_),
    .Y(_01447_));
 sky130_vsdinv _25792_ (.A(_20828_),
    .Y(_20834_));
 sky130_fd_sc_hd__a31o_1 _25793_ (.A1(_20834_),
    .A2(_20042_),
    .A3(\decoded_imm[24] ),
    .B1(_20829_),
    .X(_20835_));
 sky130_fd_sc_hd__nor2_1 _25794_ (.A(_20039_),
    .B(\decoded_imm[26] ),
    .Y(_20836_));
 sky130_fd_sc_hd__nor2_1 _25795_ (.A(_20509_),
    .B(_20663_),
    .Y(_20837_));
 sky130_fd_sc_hd__nor2_1 _25796_ (.A(_20836_),
    .B(_20837_),
    .Y(_20838_));
 sky130_fd_sc_hd__nand2_1 _25797_ (.A(_20831_),
    .B(_20822_),
    .Y(_20839_));
 sky130_fd_sc_hd__a21oi_4 _25798_ (.A1(_20819_),
    .A2(_20823_),
    .B1(_20839_),
    .Y(_20840_));
 sky130_fd_sc_hd__or3_2 _25799_ (.A(_20835_),
    .B(_20838_),
    .C(_20840_),
    .X(_20841_));
 sky130_fd_sc_hd__o21ai_1 _25800_ (.A1(_20835_),
    .A2(_20840_),
    .B1(_20838_),
    .Y(_20842_));
 sky130_fd_sc_hd__and2_1 _25801_ (.A(_20841_),
    .B(_20842_),
    .X(_01449_));
 sky130_vsdinv _25802_ (.A(\reg_pc[27] ),
    .Y(_20843_));
 sky130_fd_sc_hd__nor2_1 _25803_ (.A(_20820_),
    .B(_20843_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _25804_ (.A(net325),
    .B(\decoded_imm[27] ),
    .Y(_20844_));
 sky130_fd_sc_hd__nor2_1 _25805_ (.A(_20522_),
    .B(_20664_),
    .Y(_20845_));
 sky130_fd_sc_hd__nor2_2 _25806_ (.A(_20844_),
    .B(_20845_),
    .Y(_20846_));
 sky130_fd_sc_hd__o21ai_1 _25807_ (.A1(_20509_),
    .A2(_20663_),
    .B1(_20842_),
    .Y(_20847_));
 sky130_fd_sc_hd__xor2_1 _25808_ (.A(_20846_),
    .B(_20847_),
    .X(_01452_));
 sky130_vsdinv _25809_ (.A(\reg_pc[28] ),
    .Y(_20848_));
 sky130_fd_sc_hd__nor2_1 _25810_ (.A(_20820_),
    .B(_20848_),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _25811_ (.A(_20038_),
    .B(\decoded_imm[28] ),
    .Y(_20849_));
 sky130_fd_sc_hd__nor2_4 _25812_ (.A(_20505_),
    .B(_20665_),
    .Y(_20850_));
 sky130_fd_sc_hd__nor2_1 _25813_ (.A(_20849_),
    .B(_20850_),
    .Y(_20851_));
 sky130_fd_sc_hd__nand2_1 _25814_ (.A(_20838_),
    .B(_20846_),
    .Y(_20852_));
 sky130_fd_sc_hd__o21bai_2 _25815_ (.A1(_20835_),
    .A2(_20840_),
    .B1_N(_20852_),
    .Y(_20853_));
 sky130_vsdinv _25816_ (.A(_20845_),
    .Y(_20854_));
 sky130_fd_sc_hd__o31a_1 _25817_ (.A1(_20509_),
    .A2(_20663_),
    .A3(_20844_),
    .B1(_20854_),
    .X(_20855_));
 sky130_fd_sc_hd__nand2_1 _25818_ (.A(_20853_),
    .B(_20855_),
    .Y(_20856_));
 sky130_fd_sc_hd__xor2_1 _25819_ (.A(_20851_),
    .B(_20856_),
    .X(_01455_));
 sky130_vsdinv _25820_ (.A(\reg_pc[29] ),
    .Y(_20857_));
 sky130_fd_sc_hd__nor2_1 _25821_ (.A(_20820_),
    .B(_20857_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _25822_ (.A(_20518_),
    .B(_20666_),
    .Y(_20858_));
 sky130_fd_sc_hd__nand2_1 _25823_ (.A(_20037_),
    .B(\decoded_imm[29] ),
    .Y(_20859_));
 sky130_fd_sc_hd__nand2_1 _25824_ (.A(_20858_),
    .B(_20859_),
    .Y(_20860_));
 sky130_fd_sc_hd__a22oi_4 _25825_ (.A1(_20505_),
    .A2(_20665_),
    .B1(_20853_),
    .B2(_20855_),
    .Y(_20861_));
 sky130_fd_sc_hd__or3_2 _25826_ (.A(_20850_),
    .B(_20860_),
    .C(_20861_),
    .X(_20862_));
 sky130_fd_sc_hd__o21ai_1 _25827_ (.A1(_20850_),
    .A2(_20861_),
    .B1(_20860_),
    .Y(_20863_));
 sky130_fd_sc_hd__nand2_1 _25828_ (.A(_20862_),
    .B(_20863_),
    .Y(_01458_));
 sky130_vsdinv _25829_ (.A(\reg_pc[30] ),
    .Y(_20864_));
 sky130_fd_sc_hd__nor2_1 _25830_ (.A(_20023_),
    .B(_20864_),
    .Y(_01459_));
 sky130_fd_sc_hd__nor2_1 _25831_ (.A(_20036_),
    .B(\decoded_imm[30] ),
    .Y(_20865_));
 sky130_fd_sc_hd__nor2_2 _25832_ (.A(_20529_),
    .B(_20667_),
    .Y(_20866_));
 sky130_fd_sc_hd__nor2_1 _25833_ (.A(_20865_),
    .B(_20866_),
    .Y(_20867_));
 sky130_fd_sc_hd__o22ai_4 _25834_ (.A1(_20037_),
    .A2(\decoded_imm[29] ),
    .B1(_20850_),
    .B2(_20861_),
    .Y(_20868_));
 sky130_fd_sc_hd__nand2_1 _25835_ (.A(_20868_),
    .B(_20859_),
    .Y(_20869_));
 sky130_fd_sc_hd__xor2_1 _25836_ (.A(_20867_),
    .B(_20869_),
    .X(_01461_));
 sky130_vsdinv _25837_ (.A(\reg_pc[31] ),
    .Y(_20870_));
 sky130_fd_sc_hd__nor2_1 _25838_ (.A(_20023_),
    .B(_20870_),
    .Y(_01462_));
 sky130_fd_sc_hd__a22oi_1 _25839_ (.A1(_20529_),
    .A2(_20667_),
    .B1(_20868_),
    .B2(_20859_),
    .Y(_20871_));
 sky130_fd_sc_hd__xnor2_1 _25840_ (.A(net330),
    .B(\decoded_imm[31] ),
    .Y(_20872_));
 sky130_vsdinv _25841_ (.A(_20872_),
    .Y(_20873_));
 sky130_fd_sc_hd__o21bai_1 _25842_ (.A1(_20866_),
    .A2(_20871_),
    .B1_N(_20873_),
    .Y(_20874_));
 sky130_fd_sc_hd__a21o_1 _25843_ (.A1(_20868_),
    .A2(_20859_),
    .B1(_20865_),
    .X(_20875_));
 sky130_fd_sc_hd__nor2_1 _25844_ (.A(_20866_),
    .B(_20872_),
    .Y(_20876_));
 sky130_fd_sc_hd__nand2_1 _25845_ (.A(_20875_),
    .B(_20876_),
    .Y(_20877_));
 sky130_fd_sc_hd__nand2_1 _25846_ (.A(_20874_),
    .B(_20877_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_1 _25847_ (.A(_20555_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and2_1 _25848_ (.A(_20555_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__buf_2 _25849_ (.A(_18761_),
    .X(_20878_));
 sky130_fd_sc_hd__a21oi_1 _25850_ (.A1(_20555_),
    .A2(_01473_),
    .B1(_20878_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_1 _25851_ (.A(_20555_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__clkbuf_2 _25852_ (.A(_20554_),
    .X(_20879_));
 sky130_fd_sc_hd__and2_1 _25853_ (.A(_20879_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__and2_1 _25854_ (.A(_20879_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__and2_1 _25855_ (.A(_20879_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__and2_1 _25856_ (.A(_20879_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_1 _25857_ (.A(_20879_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_1 _25858_ (.A(_20879_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_2 _25859_ (.A(_20554_),
    .X(_20880_));
 sky130_fd_sc_hd__and2_1 _25860_ (.A(_20880_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__and2_1 _25861_ (.A(_20880_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_1 _25862_ (.A(_20880_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_1 _25863_ (.A(_20880_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__and2_1 _25864_ (.A(_20880_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_1 _25865_ (.A(_20880_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__clkbuf_2 _25866_ (.A(_20554_),
    .X(_20881_));
 sky130_fd_sc_hd__and2_1 _25867_ (.A(_20881_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_1 _25868_ (.A(_20881_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_1 _25869_ (.A(_20881_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__and2_1 _25870_ (.A(_20881_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_1 _25871_ (.A(_20881_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_1 _25872_ (.A(_20881_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__clkbuf_2 _25873_ (.A(latched_branch),
    .X(_20882_));
 sky130_fd_sc_hd__and2_1 _25874_ (.A(_20882_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__and2_1 _25875_ (.A(_20882_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_1 _25876_ (.A(_20882_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_1 _25877_ (.A(_20882_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and2_1 _25878_ (.A(_20882_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_1 _25879_ (.A(_20882_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_1 _25880_ (.A(_20554_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_1 _25881_ (.A(_20554_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__or2_1 _25882_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .X(_20883_));
 sky130_fd_sc_hd__nand2_1 _25883_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .Y(_20884_));
 sky130_fd_sc_hd__and2_1 _25884_ (.A(_20883_),
    .B(_20884_),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _25885_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .Y(_20885_));
 sky130_fd_sc_hd__and2_1 _25886_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .X(_20886_));
 sky130_fd_sc_hd__nor2_1 _25887_ (.A(_20885_),
    .B(_20886_),
    .Y(_20887_));
 sky130_fd_sc_hd__xnor2_1 _25888_ (.A(_20884_),
    .B(_20887_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _25889_ (.A(_01561_),
    .B(_02410_),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_1 _25890_ (.A(_02571_),
    .B(_02560_),
    .Y(_20888_));
 sky130_fd_sc_hd__nand2_1 _25891_ (.A(_02571_),
    .B(_02560_),
    .Y(_20889_));
 sky130_vsdinv _25892_ (.A(_20889_),
    .Y(_20890_));
 sky130_fd_sc_hd__nor2_1 _25893_ (.A(_20888_),
    .B(_20890_),
    .Y(_01567_));
 sky130_fd_sc_hd__xor2_1 _25894_ (.A(_02571_),
    .B(\decoded_imm_uj[3] ),
    .X(_20891_));
 sky130_fd_sc_hd__a31o_1 _25895_ (.A1(_20887_),
    .A2(_02590_),
    .A3(\decoded_imm_uj[1] ),
    .B1(_20886_),
    .X(_20892_));
 sky130_fd_sc_hd__xor2_1 _25896_ (.A(_20891_),
    .B(_20892_),
    .X(_01568_));
 sky130_fd_sc_hd__nor2_2 _25897_ (.A(_01475_),
    .B(_20889_),
    .Y(_20893_));
 sky130_fd_sc_hd__nor2_1 _25898_ (.A(_02582_),
    .B(_20890_),
    .Y(_20894_));
 sky130_fd_sc_hd__nor2_1 _25899_ (.A(_20893_),
    .B(_20894_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_2 _25900_ (.A(_01475_),
    .B(_00367_),
    .Y(_20895_));
 sky130_fd_sc_hd__nor2_1 _25901_ (.A(\decoded_imm_uj[4] ),
    .B(_02582_),
    .Y(_20896_));
 sky130_fd_sc_hd__or2_1 _25902_ (.A(_20895_),
    .B(_20896_),
    .X(_20897_));
 sky130_fd_sc_hd__o21a_1 _25903_ (.A1(_02571_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_20892_),
    .X(_20898_));
 sky130_fd_sc_hd__a21oi_2 _25904_ (.A1(_02571_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_20898_),
    .Y(_20899_));
 sky130_fd_sc_hd__xor2_1 _25905_ (.A(_20897_),
    .B(_20899_),
    .X(_01572_));
 sky130_fd_sc_hd__nor2_1 _25906_ (.A(_02583_),
    .B(_20893_),
    .Y(_20900_));
 sky130_fd_sc_hd__and2_1 _25907_ (.A(_20893_),
    .B(_02583_),
    .X(_20901_));
 sky130_fd_sc_hd__nor2_1 _25908_ (.A(_20900_),
    .B(_20901_),
    .Y(_01575_));
 sky130_fd_sc_hd__nor2_1 _25909_ (.A(_20896_),
    .B(_20899_),
    .Y(_20902_));
 sky130_fd_sc_hd__nor2_1 _25910_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_20903_));
 sky130_fd_sc_hd__nand2_1 _25911_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_20904_));
 sky130_fd_sc_hd__or2b_1 _25912_ (.A(_20903_),
    .B_N(_20904_),
    .X(_20905_));
 sky130_fd_sc_hd__o21ai_1 _25913_ (.A1(_20895_),
    .A2(_20902_),
    .B1(_20905_),
    .Y(_20906_));
 sky130_fd_sc_hd__or3_2 _25914_ (.A(_20895_),
    .B(_20905_),
    .C(_20902_),
    .X(_20907_));
 sky130_fd_sc_hd__nand2_1 _25915_ (.A(_20906_),
    .B(_20907_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _25916_ (.A(_02584_),
    .B(_20901_),
    .Y(_20908_));
 sky130_fd_sc_hd__nand2_1 _25917_ (.A(_20901_),
    .B(_02584_),
    .Y(_20909_));
 sky130_vsdinv _25918_ (.A(_20909_),
    .Y(_20910_));
 sky130_fd_sc_hd__nor2_1 _25919_ (.A(_20908_),
    .B(_20910_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _25920_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_20911_));
 sky130_fd_sc_hd__and2_1 _25921_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .X(_20912_));
 sky130_fd_sc_hd__nor2_1 _25922_ (.A(_20911_),
    .B(_20912_),
    .Y(_20913_));
 sky130_fd_sc_hd__o21bai_1 _25923_ (.A1(_20895_),
    .A2(_20902_),
    .B1_N(_20903_),
    .Y(_20914_));
 sky130_fd_sc_hd__nand2_1 _25924_ (.A(_20914_),
    .B(_20904_),
    .Y(_20915_));
 sky130_fd_sc_hd__xor2_1 _25925_ (.A(_20913_),
    .B(_20915_),
    .X(_01580_));
 sky130_fd_sc_hd__nor2_1 _25926_ (.A(_19080_),
    .B(_20909_),
    .Y(_20916_));
 sky130_fd_sc_hd__nor2_1 _25927_ (.A(_02585_),
    .B(_20910_),
    .Y(_20917_));
 sky130_fd_sc_hd__nor2_1 _25928_ (.A(_20916_),
    .B(_20917_),
    .Y(_01583_));
 sky130_fd_sc_hd__or2_1 _25929_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .X(_20918_));
 sky130_fd_sc_hd__nand2_2 _25930_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .Y(_20919_));
 sky130_fd_sc_hd__nand2_1 _25931_ (.A(_20918_),
    .B(_20919_),
    .Y(_20920_));
 sky130_fd_sc_hd__a21oi_2 _25932_ (.A1(_20914_),
    .A2(_20904_),
    .B1(_20911_),
    .Y(_20921_));
 sky130_fd_sc_hd__nor2_1 _25933_ (.A(_20912_),
    .B(_20921_),
    .Y(_20922_));
 sky130_fd_sc_hd__xor2_1 _25934_ (.A(_20920_),
    .B(_20922_),
    .X(_01584_));
 sky130_fd_sc_hd__or2_1 _25935_ (.A(_02586_),
    .B(_20916_),
    .X(_20923_));
 sky130_fd_sc_hd__nand2_1 _25936_ (.A(_20916_),
    .B(_02586_),
    .Y(_20924_));
 sky130_fd_sc_hd__and2_1 _25937_ (.A(_20923_),
    .B(_20924_),
    .X(_01587_));
 sky130_fd_sc_hd__nor2_2 _25938_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .Y(_20925_));
 sky130_fd_sc_hd__and2_1 _25939_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .X(_20926_));
 sky130_fd_sc_hd__nor2_1 _25940_ (.A(_20925_),
    .B(_20926_),
    .Y(_20927_));
 sky130_fd_sc_hd__o21ai_2 _25941_ (.A1(_20912_),
    .A2(_20921_),
    .B1(_20918_),
    .Y(_20928_));
 sky130_fd_sc_hd__nand2_1 _25942_ (.A(_20928_),
    .B(_20919_),
    .Y(_20929_));
 sky130_fd_sc_hd__xor2_1 _25943_ (.A(_20927_),
    .B(_20929_),
    .X(_01588_));
 sky130_fd_sc_hd__nor2_2 _25944_ (.A(_19073_),
    .B(_20924_),
    .Y(_20930_));
 sky130_fd_sc_hd__and2_1 _25945_ (.A(_20924_),
    .B(_19073_),
    .X(_20931_));
 sky130_fd_sc_hd__nor2_1 _25946_ (.A(_20930_),
    .B(_20931_),
    .Y(_01591_));
 sky130_fd_sc_hd__or2_1 _25947_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .X(_20932_));
 sky130_fd_sc_hd__nand2_2 _25948_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .Y(_20933_));
 sky130_fd_sc_hd__nand2_1 _25949_ (.A(_20932_),
    .B(_20933_),
    .Y(_20934_));
 sky130_fd_sc_hd__a21oi_4 _25950_ (.A1(_20928_),
    .A2(_20919_),
    .B1(_20925_),
    .Y(_20935_));
 sky130_fd_sc_hd__nor2_1 _25951_ (.A(_20926_),
    .B(_20935_),
    .Y(_20936_));
 sky130_fd_sc_hd__xor2_1 _25952_ (.A(_20934_),
    .B(_20936_),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_1 _25953_ (.A(_02588_),
    .B(_20930_),
    .Y(_20937_));
 sky130_fd_sc_hd__and2_1 _25954_ (.A(_20930_),
    .B(_02588_),
    .X(_20938_));
 sky130_fd_sc_hd__nor2_1 _25955_ (.A(_20937_),
    .B(_20938_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_2 _25956_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .Y(_20939_));
 sky130_fd_sc_hd__and2_1 _25957_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .X(_20940_));
 sky130_fd_sc_hd__nor2_1 _25958_ (.A(_20939_),
    .B(_20940_),
    .Y(_20941_));
 sky130_fd_sc_hd__o22ai_4 _25959_ (.A1(_02587_),
    .A2(\decoded_imm_uj[9] ),
    .B1(_20926_),
    .B2(_20935_),
    .Y(_20942_));
 sky130_fd_sc_hd__nand2_1 _25960_ (.A(_20942_),
    .B(_20933_),
    .Y(_20943_));
 sky130_fd_sc_hd__xor2_1 _25961_ (.A(_20941_),
    .B(_20943_),
    .X(_01596_));
 sky130_fd_sc_hd__or2_1 _25962_ (.A(_02589_),
    .B(_20938_),
    .X(_20944_));
 sky130_fd_sc_hd__nand2_1 _25963_ (.A(_20938_),
    .B(_02589_),
    .Y(_20945_));
 sky130_fd_sc_hd__and2_1 _25964_ (.A(_20944_),
    .B(_20945_),
    .X(_01599_));
 sky130_vsdinv _25965_ (.A(\decoded_imm_uj[11] ),
    .Y(_20946_));
 sky130_fd_sc_hd__nor2_2 _25966_ (.A(_02589_),
    .B(_20946_),
    .Y(_20947_));
 sky130_fd_sc_hd__nor2_2 _25967_ (.A(\decoded_imm_uj[11] ),
    .B(_19069_),
    .Y(_20948_));
 sky130_fd_sc_hd__a21oi_4 _25968_ (.A1(_20942_),
    .A2(_20933_),
    .B1(_20939_),
    .Y(_20949_));
 sky130_fd_sc_hd__or4_1 _25969_ (.A(_20940_),
    .B(_20947_),
    .C(_20948_),
    .D(_20949_),
    .X(_20950_));
 sky130_fd_sc_hd__o22ai_4 _25970_ (.A1(_20947_),
    .A2(_20948_),
    .B1(_20940_),
    .B2(_20949_),
    .Y(_20951_));
 sky130_fd_sc_hd__and2_1 _25971_ (.A(_20950_),
    .B(_20951_),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_2 _25972_ (.A(_19067_),
    .B(_20945_),
    .Y(_20952_));
 sky130_fd_sc_hd__and2_1 _25973_ (.A(_20945_),
    .B(_19067_),
    .X(_20953_));
 sky130_fd_sc_hd__nor2_1 _25974_ (.A(_20952_),
    .B(_20953_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _25975_ (.A(_19069_),
    .B(_20946_),
    .Y(_20954_));
 sky130_vsdinv _25976_ (.A(_20954_),
    .Y(_20955_));
 sky130_fd_sc_hd__nor2_1 _25977_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .Y(_20956_));
 sky130_fd_sc_hd__and2_1 _25978_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .X(_20957_));
 sky130_fd_sc_hd__or2_2 _25979_ (.A(_20956_),
    .B(_20957_),
    .X(_20958_));
 sky130_fd_sc_hd__a21oi_4 _25980_ (.A1(_20951_),
    .A2(_20955_),
    .B1(_20958_),
    .Y(_20959_));
 sky130_fd_sc_hd__and3_1 _25981_ (.A(_20951_),
    .B(_20955_),
    .C(_20958_),
    .X(_20960_));
 sky130_fd_sc_hd__nor2_1 _25982_ (.A(_20959_),
    .B(_20960_),
    .Y(_01604_));
 sky130_fd_sc_hd__or2_1 _25983_ (.A(_02562_),
    .B(_20952_),
    .X(_20961_));
 sky130_fd_sc_hd__nand2_2 _25984_ (.A(_20952_),
    .B(_02562_),
    .Y(_20962_));
 sky130_fd_sc_hd__and2_1 _25985_ (.A(_20961_),
    .B(_20962_),
    .X(_01607_));
 sky130_vsdinv _25986_ (.A(\decoded_imm_uj[13] ),
    .Y(_20963_));
 sky130_fd_sc_hd__nor2_2 _25987_ (.A(_02562_),
    .B(_20963_),
    .Y(_20964_));
 sky130_fd_sc_hd__nor2_2 _25988_ (.A(\decoded_imm_uj[13] ),
    .B(_19065_),
    .Y(_20965_));
 sky130_fd_sc_hd__or4_1 _25989_ (.A(_20957_),
    .B(_20964_),
    .C(_20965_),
    .D(_20959_),
    .X(_20966_));
 sky130_fd_sc_hd__o22ai_4 _25990_ (.A1(_20964_),
    .A2(_20965_),
    .B1(_20957_),
    .B2(_20959_),
    .Y(_20967_));
 sky130_fd_sc_hd__and2_1 _25991_ (.A(_20966_),
    .B(_20967_),
    .X(_01608_));
 sky130_fd_sc_hd__nor2_4 _25992_ (.A(_19061_),
    .B(_20962_),
    .Y(_20968_));
 sky130_fd_sc_hd__and2_1 _25993_ (.A(_20962_),
    .B(_19061_),
    .X(_20969_));
 sky130_fd_sc_hd__nor2_1 _25994_ (.A(_20968_),
    .B(_20969_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _25995_ (.A(_19065_),
    .B(_20963_),
    .Y(_20970_));
 sky130_vsdinv _25996_ (.A(_20970_),
    .Y(_20971_));
 sky130_fd_sc_hd__nor2_1 _25997_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .Y(_20972_));
 sky130_fd_sc_hd__and2_2 _25998_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .X(_20973_));
 sky130_fd_sc_hd__or2_2 _25999_ (.A(_20972_),
    .B(_20973_),
    .X(_20974_));
 sky130_fd_sc_hd__a21oi_4 _26000_ (.A1(_20967_),
    .A2(_20971_),
    .B1(_20974_),
    .Y(_20975_));
 sky130_fd_sc_hd__and3_1 _26001_ (.A(_20967_),
    .B(_20971_),
    .C(_20974_),
    .X(_20976_));
 sky130_fd_sc_hd__nor2_1 _26002_ (.A(_20975_),
    .B(_20976_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _26003_ (.A(_02564_),
    .B(_20968_),
    .Y(_20977_));
 sky130_fd_sc_hd__nand2_1 _26004_ (.A(_20968_),
    .B(_02564_),
    .Y(_20978_));
 sky130_vsdinv _26005_ (.A(_20978_),
    .Y(_20979_));
 sky130_fd_sc_hd__nor2_1 _26006_ (.A(_20977_),
    .B(_20979_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_2 _26007_ (.A(_02564_),
    .B(_19966_),
    .Y(_20980_));
 sky130_fd_sc_hd__nor2_2 _26008_ (.A(\decoded_imm_uj[15] ),
    .B(_19058_),
    .Y(_20981_));
 sky130_fd_sc_hd__or4_1 _26009_ (.A(_20973_),
    .B(_20980_),
    .C(_20981_),
    .D(_20975_),
    .X(_20982_));
 sky130_fd_sc_hd__o22ai_4 _26010_ (.A1(_20980_),
    .A2(_20981_),
    .B1(_20973_),
    .B2(_20975_),
    .Y(_20983_));
 sky130_fd_sc_hd__and2_1 _26011_ (.A(_20982_),
    .B(_20983_),
    .X(_01616_));
 sky130_fd_sc_hd__nor2_2 _26012_ (.A(_19056_),
    .B(_20978_),
    .Y(_20984_));
 sky130_fd_sc_hd__nor2_1 _26013_ (.A(_02565_),
    .B(_20979_),
    .Y(_20985_));
 sky130_fd_sc_hd__nor2_1 _26014_ (.A(_20984_),
    .B(_20985_),
    .Y(_01619_));
 sky130_fd_sc_hd__nor2_1 _26015_ (.A(_19058_),
    .B(_19966_),
    .Y(_20986_));
 sky130_vsdinv _26016_ (.A(_20986_),
    .Y(_20987_));
 sky130_fd_sc_hd__nor2_1 _26017_ (.A(_02565_),
    .B(\decoded_imm_uj[16] ),
    .Y(_20988_));
 sky130_fd_sc_hd__nor2_4 _26018_ (.A(_19056_),
    .B(_19965_),
    .Y(_20989_));
 sky130_fd_sc_hd__nor2_1 _26019_ (.A(_20988_),
    .B(_20989_),
    .Y(_20990_));
 sky130_vsdinv _26020_ (.A(_20990_),
    .Y(_20991_));
 sky130_fd_sc_hd__a21oi_4 _26021_ (.A1(_20983_),
    .A2(_20987_),
    .B1(_20991_),
    .Y(_20992_));
 sky130_fd_sc_hd__and3_1 _26022_ (.A(_20983_),
    .B(_20987_),
    .C(_20991_),
    .X(_20993_));
 sky130_fd_sc_hd__nor2_1 _26023_ (.A(_20992_),
    .B(_20993_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _26024_ (.A(_02566_),
    .B(_20984_),
    .Y(_20994_));
 sky130_fd_sc_hd__nand2_1 _26025_ (.A(_20984_),
    .B(_02566_),
    .Y(_20995_));
 sky130_vsdinv _26026_ (.A(_20995_),
    .Y(_20996_));
 sky130_fd_sc_hd__nor2_1 _26027_ (.A(_20994_),
    .B(_20996_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_2 _26028_ (.A(_02566_),
    .B(_19964_),
    .Y(_20997_));
 sky130_fd_sc_hd__nor2_2 _26029_ (.A(\decoded_imm_uj[17] ),
    .B(_19054_),
    .Y(_20998_));
 sky130_fd_sc_hd__or4_1 _26030_ (.A(_20989_),
    .B(_20997_),
    .C(_20998_),
    .D(_20992_),
    .X(_20999_));
 sky130_fd_sc_hd__o22ai_4 _26031_ (.A1(_20997_),
    .A2(_20998_),
    .B1(_20989_),
    .B2(_20992_),
    .Y(_21000_));
 sky130_fd_sc_hd__and2_1 _26032_ (.A(_20999_),
    .B(_21000_),
    .X(_01624_));
 sky130_fd_sc_hd__nor2_2 _26033_ (.A(_19052_),
    .B(_20995_),
    .Y(_21001_));
 sky130_fd_sc_hd__nor2_1 _26034_ (.A(_02567_),
    .B(_20996_),
    .Y(_21002_));
 sky130_fd_sc_hd__nor2_1 _26035_ (.A(_21001_),
    .B(_21002_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _26036_ (.A(_02567_),
    .B(\decoded_imm_uj[18] ),
    .Y(_21003_));
 sky130_fd_sc_hd__nor2_4 _26037_ (.A(_19052_),
    .B(_19963_),
    .Y(_21004_));
 sky130_fd_sc_hd__nor2_1 _26038_ (.A(_21003_),
    .B(_21004_),
    .Y(_21005_));
 sky130_fd_sc_hd__nor2_1 _26039_ (.A(_19054_),
    .B(_19964_),
    .Y(_21006_));
 sky130_vsdinv _26040_ (.A(_21006_),
    .Y(_21007_));
 sky130_fd_sc_hd__nand2_1 _26041_ (.A(_21000_),
    .B(_21007_),
    .Y(_21008_));
 sky130_fd_sc_hd__xor2_1 _26042_ (.A(_21005_),
    .B(_21008_),
    .X(_01628_));
 sky130_fd_sc_hd__nor2_1 _26043_ (.A(_02568_),
    .B(_21001_),
    .Y(_21009_));
 sky130_fd_sc_hd__nand2_1 _26044_ (.A(_21001_),
    .B(_02568_),
    .Y(_21010_));
 sky130_vsdinv _26045_ (.A(_21010_),
    .Y(_21011_));
 sky130_fd_sc_hd__nor2_1 _26046_ (.A(_21009_),
    .B(_21011_),
    .Y(_01631_));
 sky130_vsdinv _26047_ (.A(\decoded_imm_uj[19] ),
    .Y(_21012_));
 sky130_fd_sc_hd__nor2_2 _26048_ (.A(_02568_),
    .B(_21012_),
    .Y(_21013_));
 sky130_fd_sc_hd__nor2_2 _26049_ (.A(\decoded_imm_uj[19] ),
    .B(_19050_),
    .Y(_21014_));
 sky130_fd_sc_hd__a22oi_4 _26050_ (.A1(_19052_),
    .A2(_19963_),
    .B1(_21000_),
    .B2(_21007_),
    .Y(_21015_));
 sky130_fd_sc_hd__or4_1 _26051_ (.A(_21004_),
    .B(_21013_),
    .C(_21014_),
    .D(_21015_),
    .X(_21016_));
 sky130_fd_sc_hd__o22ai_4 _26052_ (.A1(_21013_),
    .A2(_21014_),
    .B1(_21004_),
    .B2(_21015_),
    .Y(_21017_));
 sky130_fd_sc_hd__and2_1 _26053_ (.A(_21016_),
    .B(_21017_),
    .X(_01632_));
 sky130_fd_sc_hd__nor2_1 _26054_ (.A(_19045_),
    .B(_21010_),
    .Y(_21018_));
 sky130_fd_sc_hd__nor2_1 _26055_ (.A(_02569_),
    .B(_21011_),
    .Y(_21019_));
 sky130_fd_sc_hd__nor2_1 _26056_ (.A(_21018_),
    .B(_21019_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _26057_ (.A(_19050_),
    .B(_21012_),
    .Y(_21020_));
 sky130_vsdinv _26058_ (.A(_21020_),
    .Y(_21021_));
 sky130_fd_sc_hd__nor2_1 _26059_ (.A(_02569_),
    .B(_19961_),
    .Y(_21022_));
 sky130_vsdinv _26060_ (.A(\decoded_imm_uj[20] ),
    .Y(_21023_));
 sky130_fd_sc_hd__clkbuf_4 _26061_ (.A(_21023_),
    .X(_21024_));
 sky130_fd_sc_hd__nor2_2 _26062_ (.A(_19045_),
    .B(_21024_),
    .Y(_21025_));
 sky130_fd_sc_hd__or2_1 _26063_ (.A(_21022_),
    .B(_21025_),
    .X(_21026_));
 sky130_fd_sc_hd__a21oi_1 _26064_ (.A1(_21017_),
    .A2(_21021_),
    .B1(_21026_),
    .Y(_21027_));
 sky130_fd_sc_hd__and3_1 _26065_ (.A(_21017_),
    .B(_21021_),
    .C(_21026_),
    .X(_21028_));
 sky130_fd_sc_hd__nor2_1 _26066_ (.A(_21027_),
    .B(_21028_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_1 _26067_ (.A(_02570_),
    .B(_21018_),
    .Y(_21029_));
 sky130_fd_sc_hd__and2_1 _26068_ (.A(_21018_),
    .B(_02570_),
    .X(_21030_));
 sky130_fd_sc_hd__nor2_1 _26069_ (.A(_21029_),
    .B(_21030_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _26070_ (.A(_02570_),
    .B(\decoded_imm_uj[20] ),
    .Y(_21031_));
 sky130_fd_sc_hd__nor2_1 _26071_ (.A(_19042_),
    .B(_21023_),
    .Y(_21032_));
 sky130_fd_sc_hd__or2_1 _26072_ (.A(_21031_),
    .B(_21032_),
    .X(_21033_));
 sky130_vsdinv _26073_ (.A(_21033_),
    .Y(_21034_));
 sky130_fd_sc_hd__a22oi_4 _26074_ (.A1(_19045_),
    .A2(_21024_),
    .B1(_21017_),
    .B2(_21021_),
    .Y(_21035_));
 sky130_fd_sc_hd__or2_1 _26075_ (.A(_21025_),
    .B(_21035_),
    .X(_21036_));
 sky130_fd_sc_hd__or2_1 _26076_ (.A(_21034_),
    .B(_21036_),
    .X(_21037_));
 sky130_fd_sc_hd__nand2_1 _26077_ (.A(_21036_),
    .B(_21034_),
    .Y(_21038_));
 sky130_fd_sc_hd__and2_1 _26078_ (.A(_21037_),
    .B(_21038_),
    .X(_01640_));
 sky130_fd_sc_hd__nor2_1 _26079_ (.A(_02572_),
    .B(_21030_),
    .Y(_21039_));
 sky130_fd_sc_hd__nand2_1 _26080_ (.A(_21030_),
    .B(_02572_),
    .Y(_21040_));
 sky130_vsdinv _26081_ (.A(_21040_),
    .Y(_21041_));
 sky130_fd_sc_hd__nor2_1 _26082_ (.A(_21039_),
    .B(_21041_),
    .Y(_01643_));
 sky130_fd_sc_hd__xnor2_2 _26083_ (.A(_02572_),
    .B(\decoded_imm_uj[20] ),
    .Y(_21042_));
 sky130_fd_sc_hd__a21oi_1 _26084_ (.A1(_21036_),
    .A2(_21034_),
    .B1(_21032_),
    .Y(_21043_));
 sky130_fd_sc_hd__xor2_1 _26085_ (.A(_21042_),
    .B(_21043_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_2 _26086_ (.A(_19038_),
    .B(_21040_),
    .Y(_21044_));
 sky130_fd_sc_hd__nor2_1 _26087_ (.A(_02573_),
    .B(_21041_),
    .Y(_21045_));
 sky130_fd_sc_hd__nor2_1 _26088_ (.A(_21044_),
    .B(_21045_),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _26089_ (.A(_21042_),
    .B(_21038_),
    .Y(_21046_));
 sky130_fd_sc_hd__nor2_1 _26090_ (.A(_19038_),
    .B(_21023_),
    .Y(_21047_));
 sky130_vsdinv _26091_ (.A(_21047_),
    .Y(_21048_));
 sky130_fd_sc_hd__nand2_1 _26092_ (.A(_19038_),
    .B(_21024_),
    .Y(_21049_));
 sky130_fd_sc_hd__o21a_1 _26093_ (.A1(_02572_),
    .A2(_02570_),
    .B1(_19961_),
    .X(_21050_));
 sky130_fd_sc_hd__a21o_1 _26094_ (.A1(_21048_),
    .A2(_21049_),
    .B1(_21050_),
    .X(_21051_));
 sky130_fd_sc_hd__nand2_1 _26095_ (.A(_21048_),
    .B(_21049_),
    .Y(_21052_));
 sky130_fd_sc_hd__o21bai_1 _26096_ (.A1(_21050_),
    .A2(_21046_),
    .B1_N(_21052_),
    .Y(_21053_));
 sky130_fd_sc_hd__o21a_1 _26097_ (.A1(_21046_),
    .A2(_21051_),
    .B1(_21053_),
    .X(_01648_));
 sky130_fd_sc_hd__nor2_1 _26098_ (.A(_02574_),
    .B(_21044_),
    .Y(_21054_));
 sky130_fd_sc_hd__nand2_1 _26099_ (.A(_21044_),
    .B(_02574_),
    .Y(_21055_));
 sky130_vsdinv _26100_ (.A(_21055_),
    .Y(_21056_));
 sky130_fd_sc_hd__nor2_1 _26101_ (.A(_21054_),
    .B(_21056_),
    .Y(_01651_));
 sky130_fd_sc_hd__xnor2_2 _26102_ (.A(_02574_),
    .B(_19960_),
    .Y(_21057_));
 sky130_fd_sc_hd__a21oi_1 _26103_ (.A1(_21053_),
    .A2(_21048_),
    .B1(_21057_),
    .Y(_21058_));
 sky130_fd_sc_hd__and3_1 _26104_ (.A(_21053_),
    .B(_21048_),
    .C(_21057_),
    .X(_21059_));
 sky130_fd_sc_hd__nor2_1 _26105_ (.A(_21058_),
    .B(_21059_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_2 _26106_ (.A(_19034_),
    .B(_21055_),
    .Y(_21060_));
 sky130_fd_sc_hd__nor2_1 _26107_ (.A(_02575_),
    .B(_21056_),
    .Y(_21061_));
 sky130_fd_sc_hd__nor2_1 _26108_ (.A(_21060_),
    .B(_21061_),
    .Y(_01655_));
 sky130_fd_sc_hd__buf_2 _26109_ (.A(_21024_),
    .X(_21062_));
 sky130_fd_sc_hd__nor2_2 _26110_ (.A(_02575_),
    .B(_21062_),
    .Y(_21063_));
 sky130_fd_sc_hd__nor2_2 _26111_ (.A(_19960_),
    .B(_19034_),
    .Y(_21064_));
 sky130_fd_sc_hd__or2_1 _26112_ (.A(_21063_),
    .B(_21064_),
    .X(_21065_));
 sky130_vsdinv _26113_ (.A(_21042_),
    .Y(_21066_));
 sky130_fd_sc_hd__nor2_2 _26114_ (.A(_21057_),
    .B(_21052_),
    .Y(_21067_));
 sky130_fd_sc_hd__o2111ai_4 _26115_ (.A1(_21025_),
    .A2(_21035_),
    .B1(_21034_),
    .C1(_21066_),
    .D1(_21067_),
    .Y(_21068_));
 sky130_fd_sc_hd__a41o_1 _26116_ (.A1(_19036_),
    .A2(_19038_),
    .A3(_19040_),
    .A4(_19042_),
    .B1(_21024_),
    .X(_21069_));
 sky130_fd_sc_hd__nand2_2 _26117_ (.A(_21068_),
    .B(_21069_),
    .Y(_21070_));
 sky130_fd_sc_hd__or2_1 _26118_ (.A(_21065_),
    .B(_21070_),
    .X(_21071_));
 sky130_fd_sc_hd__nand2_1 _26119_ (.A(_21070_),
    .B(_21065_),
    .Y(_21072_));
 sky130_fd_sc_hd__and2_1 _26120_ (.A(_21071_),
    .B(_21072_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_1 _26121_ (.A(_02576_),
    .B(_21060_),
    .Y(_21073_));
 sky130_fd_sc_hd__nand2_1 _26122_ (.A(_21060_),
    .B(_02576_),
    .Y(_21074_));
 sky130_vsdinv _26123_ (.A(_21074_),
    .Y(_21075_));
 sky130_fd_sc_hd__nor2_1 _26124_ (.A(_21073_),
    .B(_21075_),
    .Y(_01659_));
 sky130_fd_sc_hd__xor2_4 _26125_ (.A(_02576_),
    .B(_19960_),
    .X(_21076_));
 sky130_fd_sc_hd__o21ai_1 _26126_ (.A1(_19034_),
    .A2(_21062_),
    .B1(_21072_),
    .Y(_21077_));
 sky130_fd_sc_hd__xor2_1 _26127_ (.A(_21076_),
    .B(_21077_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_2 _26128_ (.A(_19027_),
    .B(_21074_),
    .Y(_21078_));
 sky130_fd_sc_hd__nor2_1 _26129_ (.A(_02577_),
    .B(_21075_),
    .Y(_21079_));
 sky130_fd_sc_hd__nor2_1 _26130_ (.A(_21078_),
    .B(_21079_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand3_2 _26131_ (.A(_21070_),
    .B(_21065_),
    .C(_21076_),
    .Y(_21080_));
 sky130_fd_sc_hd__o21ai_1 _26132_ (.A1(_02576_),
    .A2(_02575_),
    .B1(_19962_),
    .Y(_21081_));
 sky130_fd_sc_hd__nor2_1 _26133_ (.A(_02577_),
    .B(_19960_),
    .Y(_21082_));
 sky130_fd_sc_hd__nor2_1 _26134_ (.A(_19027_),
    .B(_21024_),
    .Y(_21083_));
 sky130_fd_sc_hd__or2_2 _26135_ (.A(_21082_),
    .B(_21083_),
    .X(_21084_));
 sky130_fd_sc_hd__a21oi_2 _26136_ (.A1(_21080_),
    .A2(_21081_),
    .B1(_21084_),
    .Y(_21085_));
 sky130_fd_sc_hd__and3_1 _26137_ (.A(_21080_),
    .B(_21084_),
    .C(_21081_),
    .X(_21086_));
 sky130_fd_sc_hd__nor2_1 _26138_ (.A(_21085_),
    .B(_21086_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _26139_ (.A(_02578_),
    .B(_21078_),
    .Y(_21087_));
 sky130_fd_sc_hd__nand2_1 _26140_ (.A(_21078_),
    .B(_02578_),
    .Y(_21088_));
 sky130_vsdinv _26141_ (.A(_21088_),
    .Y(_21089_));
 sky130_fd_sc_hd__nor2_1 _26142_ (.A(_21087_),
    .B(_21089_),
    .Y(_01667_));
 sky130_fd_sc_hd__xnor2_2 _26143_ (.A(_02578_),
    .B(_19960_),
    .Y(_21090_));
 sky130_fd_sc_hd__a211o_1 _26144_ (.A1(_02577_),
    .A2(_19962_),
    .B1(_21090_),
    .C1(_21085_),
    .X(_21091_));
 sky130_fd_sc_hd__o21ai_1 _26145_ (.A1(_21083_),
    .A2(_21085_),
    .B1(_21090_),
    .Y(_21092_));
 sky130_fd_sc_hd__nand2_1 _26146_ (.A(_21091_),
    .B(_21092_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _26147_ (.A(_19023_),
    .B(_21088_),
    .Y(_21093_));
 sky130_fd_sc_hd__nor2_1 _26148_ (.A(_02579_),
    .B(_21089_),
    .Y(_21094_));
 sky130_fd_sc_hd__nor2_1 _26149_ (.A(_21093_),
    .B(_21094_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _26150_ (.A(_02579_),
    .B(_19961_),
    .Y(_21095_));
 sky130_fd_sc_hd__nor2_1 _26151_ (.A(_19023_),
    .B(_21062_),
    .Y(_21096_));
 sky130_fd_sc_hd__or2_1 _26152_ (.A(_21095_),
    .B(_21096_),
    .X(_21097_));
 sky130_vsdinv _26153_ (.A(_21097_),
    .Y(_21098_));
 sky130_fd_sc_hd__nor2_2 _26154_ (.A(_21090_),
    .B(_21084_),
    .Y(_21099_));
 sky130_fd_sc_hd__o2111ai_4 _26155_ (.A1(_21063_),
    .A2(_21064_),
    .B1(_21076_),
    .C1(_21099_),
    .D1(_21070_),
    .Y(_21100_));
 sky130_fd_sc_hd__a41o_1 _26156_ (.A1(_19025_),
    .A2(_19027_),
    .A3(_19030_),
    .A4(_19034_),
    .B1(_21062_),
    .X(_21101_));
 sky130_fd_sc_hd__nand2_2 _26157_ (.A(_21100_),
    .B(_21101_),
    .Y(_21102_));
 sky130_fd_sc_hd__nor2_1 _26158_ (.A(_21098_),
    .B(_21102_),
    .Y(_04073_));
 sky130_fd_sc_hd__nand2_1 _26159_ (.A(_21102_),
    .B(_21098_),
    .Y(_04074_));
 sky130_fd_sc_hd__nor2b_1 _26160_ (.A(_04073_),
    .B_N(_04074_),
    .Y(_01672_));
 sky130_fd_sc_hd__or2_1 _26161_ (.A(_02580_),
    .B(_21093_),
    .X(_04075_));
 sky130_fd_sc_hd__nand2_1 _26162_ (.A(_21093_),
    .B(_02580_),
    .Y(_04076_));
 sky130_fd_sc_hd__and2_1 _26163_ (.A(_04075_),
    .B(_04076_),
    .X(_01675_));
 sky130_vsdinv _26164_ (.A(_21096_),
    .Y(_04077_));
 sky130_fd_sc_hd__nor2_2 _26165_ (.A(_02580_),
    .B(_19961_),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _26166_ (.A(_19021_),
    .B(_21062_),
    .Y(_04079_));
 sky130_fd_sc_hd__o2bb2ai_1 _26167_ (.A1_N(_04077_),
    .A2_N(_04074_),
    .B1(_04078_),
    .B2(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__nor2_1 _26168_ (.A(_04078_),
    .B(_04079_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand3_1 _26169_ (.A(_04074_),
    .B(_04077_),
    .C(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _26170_ (.A(_04080_),
    .B(_04082_),
    .Y(_01676_));
 sky130_fd_sc_hd__xor2_1 _26171_ (.A(_19018_),
    .B(_04076_),
    .X(_01679_));
 sky130_fd_sc_hd__nor2_2 _26172_ (.A(_04078_),
    .B(_21097_),
    .Y(_04083_));
 sky130_fd_sc_hd__o21a_1 _26173_ (.A1(_02580_),
    .A2(_02579_),
    .B1(_19962_),
    .X(_04084_));
 sky130_fd_sc_hd__nand2_1 _26174_ (.A(_21062_),
    .B(_02581_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _26175_ (.A(_19018_),
    .B(_19962_),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_1 _26176_ (.A(_04085_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__a211oi_2 _26177_ (.A1(_21102_),
    .A2(_04083_),
    .B1(_04084_),
    .C1(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _26178_ (.A(_21102_),
    .B(_04083_),
    .Y(_04089_));
 sky130_vsdinv _26179_ (.A(_04084_),
    .Y(_04090_));
 sky130_fd_sc_hd__a22oi_1 _26180_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_04089_),
    .B2(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__nor2_1 _26181_ (.A(_04088_),
    .B(_04091_),
    .Y(_01680_));
 sky130_fd_sc_hd__nor2_4 _26182_ (.A(\mem_wordsize[2] ),
    .B(\mem_wordsize[1] ),
    .Y(_04092_));
 sky130_fd_sc_hd__clkbuf_4 _26183_ (.A(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__buf_4 _26184_ (.A(_04093_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_2 _26185_ (.A(\mem_wordsize[2] ),
    .X(_04094_));
 sky130_fd_sc_hd__a211o_4 _26186_ (.A1(_20494_),
    .A2(_04094_),
    .B1(_00304_),
    .C1(_04093_),
    .X(net233));
 sky130_fd_sc_hd__and3_1 _26187_ (.A(net233),
    .B(_18855_),
    .C(_18853_),
    .X(_01684_));
 sky130_fd_sc_hd__and3_1 _26188_ (.A(_00301_),
    .B(_20551_),
    .C(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_4 _26189_ (.A(_20063_),
    .B(_20323_),
    .Y(_04095_));
 sky130_fd_sc_hd__a211o_4 _26190_ (.A1(_20494_),
    .A2(_04094_),
    .B1(_04092_),
    .C1(_04095_),
    .X(net234));
 sky130_fd_sc_hd__and3_1 _26191_ (.A(net234),
    .B(_18853_),
    .C(_18855_),
    .X(_01687_));
 sky130_fd_sc_hd__and3_1 _26192_ (.A(_00301_),
    .B(_20551_),
    .C(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__nor2_4 _26193_ (.A(_20064_),
    .B(_20494_),
    .Y(_04096_));
 sky130_fd_sc_hd__nor2_1 _26194_ (.A(_20494_),
    .B(_20336_),
    .Y(_04097_));
 sky130_fd_sc_hd__or3_4 _26195_ (.A(_04092_),
    .B(_04096_),
    .C(_04097_),
    .X(net235));
 sky130_fd_sc_hd__and3_1 _26196_ (.A(net235),
    .B(_18853_),
    .C(_18855_),
    .X(_01690_));
 sky130_fd_sc_hd__and3_1 _26197_ (.A(_00301_),
    .B(_20551_),
    .C(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__nor2_4 _26198_ (.A(_20494_),
    .B(_20323_),
    .Y(_04098_));
 sky130_fd_sc_hd__or3_4 _26199_ (.A(_04092_),
    .B(_04097_),
    .C(_04098_),
    .X(net236));
 sky130_fd_sc_hd__and2_1 _26200_ (.A(net232),
    .B(net236),
    .X(_01693_));
 sky130_fd_sc_hd__and3_1 _26201_ (.A(_00301_),
    .B(_20551_),
    .C(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_4 _26202_ (.A(\irq_pending[1] ),
    .B(net12),
    .Y(_01696_));
 sky130_fd_sc_hd__inv_2 _26203_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_1 _26204_ (.A(_18848_),
    .B(_01696_),
    .Y(_01698_));
 sky130_fd_sc_hd__or3_1 _26205_ (.A(\cpu_state[0] ),
    .B(_02542_),
    .C(_18777_),
    .X(_04099_));
 sky130_fd_sc_hd__nor2_1 _26206_ (.A(_20388_),
    .B(_04099_),
    .Y(_01700_));
 sky130_fd_sc_hd__nor2_1 _26207_ (.A(_20332_),
    .B(_01697_),
    .Y(_01701_));
 sky130_fd_sc_hd__a2bb2o_1 _26208_ (.A1_N(_18743_),
    .A2_N(_01704_),
    .B1(_01697_),
    .B2(_04099_),
    .X(_01705_));
 sky130_vsdinv _26209_ (.A(net33),
    .Y(_01707_));
 sky130_fd_sc_hd__clkbuf_2 _26210_ (.A(_04095_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_2 _26211_ (.A(_04096_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_2 _26212_ (.A(_04098_),
    .X(_04102_));
 sky130_fd_sc_hd__a22o_1 _26213_ (.A1(_04101_),
    .A2(net40),
    .B1(_04102_),
    .B2(net49),
    .X(_04103_));
 sky130_fd_sc_hd__a21oi_1 _26214_ (.A1(net63),
    .A2(_04100_),
    .B1(_04103_),
    .Y(_01708_));
 sky130_fd_sc_hd__clkbuf_2 _26215_ (.A(_04094_),
    .X(_04104_));
 sky130_fd_sc_hd__o2bb2a_1 _26216_ (.A1_N(_04104_),
    .A2_N(_01710_),
    .B1(_01709_),
    .B2(_20550_),
    .X(_01711_));
 sky130_vsdinv _26217_ (.A(_20005_),
    .Y(_04105_));
 sky130_fd_sc_hd__buf_2 _26218_ (.A(_04105_),
    .X(_04106_));
 sky130_vsdinv _26219_ (.A(_20009_),
    .Y(_04107_));
 sky130_fd_sc_hd__buf_2 _26220_ (.A(_04107_),
    .X(_04108_));
 sky130_vsdinv _26221_ (.A(instr_rdcycleh),
    .Y(_04109_));
 sky130_fd_sc_hd__clkbuf_2 _26222_ (.A(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__and3_4 _26223_ (.A(_04106_),
    .B(_04108_),
    .C(_04110_),
    .X(_01714_));
 sky130_fd_sc_hd__buf_2 _26224_ (.A(_04107_),
    .X(_04111_));
 sky130_fd_sc_hd__nand2_1 _26225_ (.A(\count_instr[32] ),
    .B(_20006_),
    .Y(_04112_));
 sky130_fd_sc_hd__o221a_1 _26226_ (.A1(_19111_),
    .A2(_04111_),
    .B1(_04110_),
    .B2(_19539_),
    .C1(_04112_),
    .X(_01715_));
 sky130_vsdinv _26227_ (.A(\irq_mask[0] ),
    .Y(_04113_));
 sky130_fd_sc_hd__clkbuf_2 _26228_ (.A(_18714_),
    .X(_04114_));
 sky130_fd_sc_hd__nand2_1 _26229_ (.A(_19975_),
    .B(\timer[0] ),
    .Y(_04115_));
 sky130_fd_sc_hd__o221a_1 _26230_ (.A1(_04113_),
    .A2(_04114_),
    .B1(_18709_),
    .B2(_18851_),
    .C1(_04115_),
    .X(_01718_));
 sky130_fd_sc_hd__clkbuf_4 _26231_ (.A(_18697_),
    .X(_04116_));
 sky130_fd_sc_hd__nand2_1 _26232_ (.A(_20670_),
    .B(_20669_),
    .Y(_04117_));
 sky130_fd_sc_hd__nand2_2 _26233_ (.A(\decoded_imm[0] ),
    .B(\reg_next_pc[0] ),
    .Y(_04118_));
 sky130_fd_sc_hd__clkbuf_2 _26234_ (.A(_18722_),
    .X(_04119_));
 sky130_fd_sc_hd__buf_4 _26235_ (.A(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__nor2_1 _26236_ (.A(_01712_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__clkbuf_2 _26237_ (.A(_18718_),
    .X(_04122_));
 sky130_fd_sc_hd__a2bb2o_1 _26238_ (.A1_N(_01719_),
    .A2_N(_19360_),
    .B1(_04122_),
    .B2(_01713_),
    .X(_04123_));
 sky130_fd_sc_hd__a311o_1 _26239_ (.A1(_04116_),
    .A2(_04117_),
    .A3(_04118_),
    .B1(_04121_),
    .C1(_04123_),
    .X(_01720_));
 sky130_vsdinv _26240_ (.A(net525),
    .Y(_01721_));
 sky130_fd_sc_hd__a22o_1 _26241_ (.A1(_04101_),
    .A2(net41),
    .B1(_04102_),
    .B2(net50),
    .X(_04124_));
 sky130_fd_sc_hd__a21oi_1 _26242_ (.A1(net64),
    .A2(_04100_),
    .B1(_04124_),
    .Y(_01722_));
 sky130_fd_sc_hd__o2bb2a_1 _26243_ (.A1_N(_04104_),
    .A2_N(_01724_),
    .B1(_01723_),
    .B2(_20550_),
    .X(_01725_));
 sky130_fd_sc_hd__nand2_1 _26244_ (.A(\count_instr[33] ),
    .B(_20006_),
    .Y(_04125_));
 sky130_fd_sc_hd__o221a_1 _26245_ (.A1(_19110_),
    .A2(_04111_),
    .B1(_04110_),
    .B2(_19419_),
    .C1(_04125_),
    .X(_01729_));
 sky130_fd_sc_hd__clkbuf_2 _26246_ (.A(_18712_),
    .X(_04126_));
 sky130_vsdinv _26247_ (.A(\timer[1] ),
    .Y(_04127_));
 sky130_fd_sc_hd__clkbuf_2 _26248_ (.A(_18710_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_2 _26249_ (.A(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__nand2_1 _26250_ (.A(\cpuregs_rs1[1] ),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__o221a_1 _26251_ (.A1(_18848_),
    .A2(_04114_),
    .B1(_04126_),
    .B2(_04127_),
    .C1(_04130_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_1 _26252_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _26253_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04132_));
 sky130_fd_sc_hd__or2b_1 _26254_ (.A(_04131_),
    .B_N(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__or2_1 _26255_ (.A(_04118_),
    .B(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__nand2_1 _26256_ (.A(_04133_),
    .B(_04118_),
    .Y(_04135_));
 sky130_fd_sc_hd__buf_2 _26257_ (.A(_20387_),
    .X(_04136_));
 sky130_fd_sc_hd__o22a_1 _26258_ (.A1(_01726_),
    .A2(_04119_),
    .B1(_19335_),
    .B2(_01732_),
    .X(_04137_));
 sky130_fd_sc_hd__a21bo_1 _26259_ (.A1(_04136_),
    .A2(_01727_),
    .B1_N(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__a31o_1 _26260_ (.A1(_04134_),
    .A2(_20390_),
    .A3(_04135_),
    .B1(_04138_),
    .X(_01733_));
 sky130_vsdinv _26261_ (.A(net55),
    .Y(_01734_));
 sky130_fd_sc_hd__a22o_1 _26262_ (.A1(_04101_),
    .A2(net42),
    .B1(_04102_),
    .B2(net51),
    .X(_04139_));
 sky130_fd_sc_hd__a21oi_1 _26263_ (.A1(net34),
    .A2(_04100_),
    .B1(_04139_),
    .Y(_01735_));
 sky130_fd_sc_hd__o2bb2a_1 _26264_ (.A1_N(_04104_),
    .A2_N(_01737_),
    .B1(_01736_),
    .B2(_20550_),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_1 _26265_ (.A(_20012_),
    .B(\count_cycle[34] ),
    .Y(_04140_));
 sky130_fd_sc_hd__o221a_1 _26266_ (.A1(_19233_),
    .A2(_04106_),
    .B1(_19109_),
    .B2(_04108_),
    .C1(_04140_),
    .X(_01742_));
 sky130_fd_sc_hd__clkbuf_2 _26267_ (.A(_04128_),
    .X(_04141_));
 sky130_fd_sc_hd__a22o_1 _26268_ (.A1(\irq_mask[2] ),
    .A2(_19985_),
    .B1(_19975_),
    .B2(\timer[2] ),
    .X(_04142_));
 sky130_fd_sc_hd__a21oi_1 _26269_ (.A1(\cpuregs_rs1[2] ),
    .A2(_04141_),
    .B1(_04142_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_2 _26270_ (.A(_02073_),
    .B(_20240_),
    .Y(_04143_));
 sky130_fd_sc_hd__nor2_2 _26271_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_04144_));
 sky130_fd_sc_hd__o21ai_2 _26272_ (.A1(_04118_),
    .A2(_04131_),
    .B1(_04132_),
    .Y(_04145_));
 sky130_fd_sc_hd__or3b_1 _26273_ (.A(_04143_),
    .B(_04144_),
    .C_N(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__buf_2 _26274_ (.A(\cpu_state[4] ),
    .X(_04147_));
 sky130_fd_sc_hd__o21bai_1 _26275_ (.A1(_04143_),
    .A2(_04144_),
    .B1_N(_04145_),
    .Y(_04148_));
 sky130_fd_sc_hd__clkbuf_2 _26276_ (.A(_18707_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_2 _26277_ (.A(_18718_),
    .X(_04150_));
 sky130_fd_sc_hd__a2bb2o_1 _26278_ (.A1_N(_01745_),
    .A2_N(_04149_),
    .B1(_04150_),
    .B2(_01740_),
    .X(_04151_));
 sky130_fd_sc_hd__nor2_1 _26279_ (.A(_01739_),
    .B(_20541_),
    .Y(_04152_));
 sky130_fd_sc_hd__a311o_1 _26280_ (.A1(_04146_),
    .A2(_04147_),
    .A3(_04148_),
    .B1(_04151_),
    .C1(_04152_),
    .X(_01746_));
 sky130_vsdinv _26281_ (.A(net58),
    .Y(_01747_));
 sky130_fd_sc_hd__a22o_1 _26282_ (.A1(_04101_),
    .A2(net526),
    .B1(_04102_),
    .B2(net52),
    .X(_04153_));
 sky130_fd_sc_hd__a21oi_1 _26283_ (.A1(net35),
    .A2(_04100_),
    .B1(_04153_),
    .Y(_01748_));
 sky130_fd_sc_hd__o2bb2a_1 _26284_ (.A1_N(_04104_),
    .A2_N(_01750_),
    .B1(_01749_),
    .B2(_20550_),
    .X(_01751_));
 sky130_fd_sc_hd__nand2_1 _26285_ (.A(\count_instr[35] ),
    .B(_20006_),
    .Y(_04154_));
 sky130_fd_sc_hd__o221a_1 _26286_ (.A1(_19304_),
    .A2(_04111_),
    .B1(_04110_),
    .B2(_19450_),
    .C1(_04154_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _26287_ (.A(\cpuregs_rs1[3] ),
    .B(_04129_),
    .Y(_04155_));
 sky130_fd_sc_hd__o221a_1 _26288_ (.A1(_18600_),
    .A2(_04114_),
    .B1(_04126_),
    .B2(_20561_),
    .C1(_04155_),
    .X(_01757_));
 sky130_fd_sc_hd__nor2_1 _26289_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _26290_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04157_));
 sky130_fd_sc_hd__or2b_1 _26291_ (.A(_04156_),
    .B_N(_04157_),
    .X(_04158_));
 sky130_vsdinv _26292_ (.A(_04144_),
    .Y(_04159_));
 sky130_fd_sc_hd__a21oi_2 _26293_ (.A1(_04145_),
    .A2(_04159_),
    .B1(_04143_),
    .Y(_04160_));
 sky130_fd_sc_hd__or2_1 _26294_ (.A(_04158_),
    .B(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_1 _26295_ (.A(_04160_),
    .B(_04158_),
    .Y(_04162_));
 sky130_fd_sc_hd__o22a_1 _26296_ (.A1(_01752_),
    .A2(_04119_),
    .B1(_19335_),
    .B2(_01758_),
    .X(_04163_));
 sky130_fd_sc_hd__a21bo_1 _26297_ (.A1(_04136_),
    .A2(_01753_),
    .B1_N(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__a31o_1 _26298_ (.A1(_04161_),
    .A2(_20390_),
    .A3(_04162_),
    .B1(_04164_),
    .X(_01759_));
 sky130_vsdinv _26299_ (.A(net59),
    .Y(_01760_));
 sky130_fd_sc_hd__a22o_1 _26300_ (.A1(_04101_),
    .A2(net524),
    .B1(_04102_),
    .B2(net53),
    .X(_04165_));
 sky130_fd_sc_hd__a21oi_1 _26301_ (.A1(net528),
    .A2(_04100_),
    .B1(_04165_),
    .Y(_01761_));
 sky130_fd_sc_hd__clkbuf_4 _26302_ (.A(_04094_),
    .X(_04166_));
 sky130_fd_sc_hd__o2bb2a_1 _26303_ (.A1_N(_04166_),
    .A2_N(_01763_),
    .B1(_01762_),
    .B2(_20550_),
    .X(_01764_));
 sky130_fd_sc_hd__clkbuf_2 _26304_ (.A(_20005_),
    .X(_04167_));
 sky130_fd_sc_hd__nand2_1 _26305_ (.A(\count_instr[36] ),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__o221a_1 _26306_ (.A1(_19306_),
    .A2(_04111_),
    .B1(_04110_),
    .B2(_19452_),
    .C1(_04168_),
    .X(_01768_));
 sky130_fd_sc_hd__a22o_1 _26307_ (.A1(\irq_mask[4] ),
    .A2(_19985_),
    .B1(_19975_),
    .B2(\timer[4] ),
    .X(_04169_));
 sky130_fd_sc_hd__a21oi_1 _26308_ (.A1(\cpuregs_rs1[4] ),
    .A2(_04141_),
    .B1(_04169_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _26309_ (.A(_20683_),
    .B(_20250_),
    .Y(_04170_));
 sky130_fd_sc_hd__nand2_1 _26310_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .Y(_04171_));
 sky130_fd_sc_hd__and2_1 _26311_ (.A(_04170_),
    .B(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__o21ai_1 _26312_ (.A1(_04156_),
    .A2(_04160_),
    .B1(_04157_),
    .Y(_04173_));
 sky130_fd_sc_hd__or2_1 _26313_ (.A(_04172_),
    .B(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__nand2_1 _26314_ (.A(_04173_),
    .B(_04172_),
    .Y(_04175_));
 sky130_fd_sc_hd__clkbuf_2 _26315_ (.A(_18722_),
    .X(_04176_));
 sky130_fd_sc_hd__o22a_1 _26316_ (.A1(_01765_),
    .A2(_04176_),
    .B1(_19335_),
    .B2(_01771_),
    .X(_04177_));
 sky130_fd_sc_hd__a21bo_1 _26317_ (.A1(_04136_),
    .A2(_01766_),
    .B1_N(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__a31o_1 _26318_ (.A1(_04174_),
    .A2(_20390_),
    .A3(_04175_),
    .B1(_04178_),
    .X(_01772_));
 sky130_vsdinv _26319_ (.A(net522),
    .Y(_01773_));
 sky130_fd_sc_hd__a22o_1 _26320_ (.A1(_04101_),
    .A2(net46),
    .B1(_04102_),
    .B2(net54),
    .X(_04179_));
 sky130_fd_sc_hd__a21oi_1 _26321_ (.A1(net37),
    .A2(_04100_),
    .B1(_04179_),
    .Y(_01774_));
 sky130_fd_sc_hd__o2bb2a_1 _26322_ (.A1_N(_04166_),
    .A2_N(_01776_),
    .B1(_01775_),
    .B2(_20549_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_2 _26323_ (.A(_04107_),
    .X(_04180_));
 sky130_fd_sc_hd__nand2_1 _26324_ (.A(_19220_),
    .B(_04167_),
    .Y(_04181_));
 sky130_fd_sc_hd__o221a_1 _26325_ (.A1(_19108_),
    .A2(_04180_),
    .B1(_04110_),
    .B2(_19453_),
    .C1(_04181_),
    .X(_01781_));
 sky130_fd_sc_hd__a22o_1 _26326_ (.A1(\irq_mask[5] ),
    .A2(_19985_),
    .B1(_19975_),
    .B2(\timer[5] ),
    .X(_04182_));
 sky130_fd_sc_hd__a21oi_1 _26327_ (.A1(\cpuregs_rs1[5] ),
    .A2(_04141_),
    .B1(_04182_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_1 _26328_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _26329_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_04184_));
 sky130_fd_sc_hd__and2b_1 _26330_ (.A_N(_04183_),
    .B(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__nand2_1 _26331_ (.A(_04175_),
    .B(_04171_),
    .Y(_04186_));
 sky130_fd_sc_hd__or2_1 _26332_ (.A(_04185_),
    .B(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__nand2_1 _26333_ (.A(_04186_),
    .B(_04185_),
    .Y(_04188_));
 sky130_fd_sc_hd__a2bb2o_1 _26334_ (.A1_N(_01784_),
    .A2_N(_04149_),
    .B1(_04150_),
    .B2(_01779_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_4 _26335_ (.A(_04119_),
    .X(_04190_));
 sky130_fd_sc_hd__nor2_1 _26336_ (.A(_01778_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__a311o_1 _26337_ (.A1(_04187_),
    .A2(_04147_),
    .A3(_04188_),
    .B1(_04189_),
    .C1(_04191_),
    .X(_01785_));
 sky130_vsdinv _26338_ (.A(net61),
    .Y(_01786_));
 sky130_fd_sc_hd__a22o_1 _26339_ (.A1(_04096_),
    .A2(net47),
    .B1(_04098_),
    .B2(net523),
    .X(_04192_));
 sky130_fd_sc_hd__a21oi_1 _26340_ (.A1(net38),
    .A2(_04095_),
    .B1(_04192_),
    .Y(_01787_));
 sky130_fd_sc_hd__o2bb2a_1 _26341_ (.A1_N(_04166_),
    .A2_N(_01789_),
    .B1(_01788_),
    .B2(_20549_),
    .X(_01790_));
 sky130_fd_sc_hd__clkbuf_2 _26342_ (.A(_04109_),
    .X(_04193_));
 sky130_fd_sc_hd__nand2_1 _26343_ (.A(\count_instr[38] ),
    .B(_04167_),
    .Y(_04194_));
 sky130_fd_sc_hd__o221a_1 _26344_ (.A1(_19103_),
    .A2(_04180_),
    .B1(_04193_),
    .B2(_19410_),
    .C1(_04194_),
    .X(_01794_));
 sky130_fd_sc_hd__a22o_1 _26345_ (.A1(\irq_mask[6] ),
    .A2(_19985_),
    .B1(_19975_),
    .B2(\timer[6] ),
    .X(_04195_));
 sky130_fd_sc_hd__a21oi_1 _26346_ (.A1(\cpuregs_rs1[6] ),
    .A2(_04141_),
    .B1(_04195_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand2_1 _26347_ (.A(_20695_),
    .B(_20640_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand2_1 _26348_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _26349_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__o21ai_1 _26350_ (.A1(_04171_),
    .A2(_04183_),
    .B1(_04184_),
    .Y(_04199_));
 sky130_fd_sc_hd__a31o_1 _26351_ (.A1(_04173_),
    .A2(_04172_),
    .A3(_04185_),
    .B1(_04199_),
    .X(_04200_));
 sky130_vsdinv _26352_ (.A(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_1 _26353_ (.A(_04198_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21o_1 _26354_ (.A1(_04201_),
    .A2(_04198_),
    .B1(_20539_),
    .X(_04203_));
 sky130_fd_sc_hd__buf_2 _26355_ (.A(_20387_),
    .X(_04204_));
 sky130_fd_sc_hd__buf_2 _26356_ (.A(_18707_),
    .X(_04205_));
 sky130_fd_sc_hd__o2bb2a_1 _26357_ (.A1_N(_04204_),
    .A2_N(_01792_),
    .B1(_01797_),
    .B2(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__o221ai_2 _26358_ (.A1(_20541_),
    .A2(_01791_),
    .B1(_04202_),
    .B2(_04203_),
    .C1(_04206_),
    .Y(_01798_));
 sky130_vsdinv _26359_ (.A(net62),
    .Y(_01799_));
 sky130_fd_sc_hd__a22o_1 _26360_ (.A1(_04096_),
    .A2(net48),
    .B1(_04098_),
    .B2(net57),
    .X(_04207_));
 sky130_fd_sc_hd__a21oi_1 _26361_ (.A1(net527),
    .A2(_04095_),
    .B1(_04207_),
    .Y(_01800_));
 sky130_fd_sc_hd__o2bb2a_1 _26362_ (.A1_N(_04166_),
    .A2_N(_01802_),
    .B1(_01801_),
    .B2(_20549_),
    .X(_01803_));
 sky130_fd_sc_hd__nand2_1 _26363_ (.A(\count_instr[39] ),
    .B(_04167_),
    .Y(_04208_));
 sky130_fd_sc_hd__o221a_1 _26364_ (.A1(_19102_),
    .A2(_04180_),
    .B1(_04193_),
    .B2(_19411_),
    .C1(_04208_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_1 _26365_ (.A(\cpuregs_rs1[7] ),
    .B(_04129_),
    .Y(_04209_));
 sky130_fd_sc_hd__o221a_1 _26366_ (.A1(_18840_),
    .A2(_04114_),
    .B1(_04126_),
    .B2(_20596_),
    .C1(_04209_),
    .X(_01809_));
 sky130_vsdinv _26367_ (.A(_01804_),
    .Y(_04210_));
 sky130_fd_sc_hd__nor2_1 _26368_ (.A(_20701_),
    .B(_20641_),
    .Y(_04211_));
 sky130_vsdinv _26369_ (.A(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__nor2_1 _26370_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_04213_));
 sky130_vsdinv _26371_ (.A(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__nand2_1 _26372_ (.A(_04212_),
    .B(_04214_),
    .Y(_04215_));
 sky130_vsdinv _26373_ (.A(_04215_),
    .Y(_04216_));
 sky130_vsdinv _26374_ (.A(_04197_),
    .Y(_04217_));
 sky130_fd_sc_hd__or2_1 _26375_ (.A(_04217_),
    .B(_04202_),
    .X(_04218_));
 sky130_fd_sc_hd__or2_1 _26376_ (.A(_04216_),
    .B(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__nand2_1 _26377_ (.A(_04218_),
    .B(_04216_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _26378_ (.A(_01810_),
    .B(_19316_),
    .Y(_04221_));
 sky130_fd_sc_hd__a31o_1 _26379_ (.A1(_04219_),
    .A2(\cpu_state[4] ),
    .A3(_04220_),
    .B1(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__a221o_1 _26380_ (.A1(_18544_),
    .A2(_04210_),
    .B1(_20388_),
    .B2(_01805_),
    .C1(_04222_),
    .X(_01811_));
 sky130_vsdinv _26381_ (.A(net63),
    .Y(_01812_));
 sky130_fd_sc_hd__clkbuf_2 _26382_ (.A(_04094_),
    .X(_04223_));
 sky130_fd_sc_hd__nand2_1 _26383_ (.A(_04223_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_8 _26384_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_vsdinv _26385_ (.A(latched_is_lh),
    .Y(_04224_));
 sky130_fd_sc_hd__clkbuf_2 _26386_ (.A(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__nand2_2 _26387_ (.A(_04210_),
    .B(latched_is_lb),
    .Y(_04226_));
 sky130_fd_sc_hd__clkbuf_2 _26388_ (.A(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__o21a_1 _26389_ (.A1(_04225_),
    .A2(_01815_),
    .B1(_04227_),
    .X(_01817_));
 sky130_fd_sc_hd__nand2_1 _26390_ (.A(\count_instr[8] ),
    .B(_20010_),
    .Y(_04228_));
 sky130_fd_sc_hd__o221a_1 _26391_ (.A1(_19224_),
    .A2(_04106_),
    .B1(_04193_),
    .B2(_19414_),
    .C1(_04228_),
    .X(_01821_));
 sky130_fd_sc_hd__nand2_1 _26392_ (.A(\cpuregs_rs1[8] ),
    .B(_04129_),
    .Y(_04229_));
 sky130_fd_sc_hd__o221a_1 _26393_ (.A1(_18628_),
    .A2(_04114_),
    .B1(_04126_),
    .B2(_20598_),
    .C1(_04229_),
    .X(_01823_));
 sky130_fd_sc_hd__nand2_1 _26394_ (.A(_20707_),
    .B(_20642_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_1 _26395_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _26396_ (.A(_04230_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__a21oi_1 _26397_ (.A1(_04214_),
    .A2(_04217_),
    .B1(_04211_),
    .Y(_04233_));
 sky130_vsdinv _26398_ (.A(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__and4_1 _26399_ (.A(_04200_),
    .B(_04197_),
    .C(_04196_),
    .D(_04216_),
    .X(_04235_));
 sky130_fd_sc_hd__nor2_1 _26400_ (.A(_04234_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__or2_1 _26401_ (.A(_04232_),
    .B(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _26402_ (.A(_04236_),
    .B(_04232_),
    .Y(_04238_));
 sky130_fd_sc_hd__clkbuf_2 _26403_ (.A(_18706_),
    .X(_04239_));
 sky130_fd_sc_hd__o22a_1 _26404_ (.A1(_01818_),
    .A2(_04176_),
    .B1(_04239_),
    .B2(_01824_),
    .X(_04240_));
 sky130_fd_sc_hd__a21bo_1 _26405_ (.A1(_04136_),
    .A2(_01819_),
    .B1_N(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__a31o_1 _26406_ (.A1(_04237_),
    .A2(_20390_),
    .A3(_04238_),
    .B1(_04241_),
    .X(_01825_));
 sky130_vsdinv _26407_ (.A(net64),
    .Y(_01826_));
 sky130_fd_sc_hd__nand2_1 _26408_ (.A(_04223_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o21a_1 _26409_ (.A1(_04225_),
    .A2(_01829_),
    .B1(_04227_),
    .X(_01830_));
 sky130_fd_sc_hd__nand2_1 _26410_ (.A(_20012_),
    .B(\count_cycle[41] ),
    .Y(_04242_));
 sky130_fd_sc_hd__o221a_1 _26411_ (.A1(_19223_),
    .A2(_04106_),
    .B1(_19106_),
    .B2(_04108_),
    .C1(_04242_),
    .X(_01834_));
 sky130_fd_sc_hd__clkbuf_2 _26412_ (.A(_19974_),
    .X(_04243_));
 sky130_fd_sc_hd__a22o_1 _26413_ (.A1(\irq_mask[9] ),
    .A2(_19985_),
    .B1(_04243_),
    .B2(\timer[9] ),
    .X(_04244_));
 sky130_fd_sc_hd__a21oi_1 _26414_ (.A1(\cpuregs_rs1[9] ),
    .A2(_04141_),
    .B1(_04244_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _26415_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_04245_));
 sky130_fd_sc_hd__nor2_1 _26416_ (.A(_20716_),
    .B(_20643_),
    .Y(_04246_));
 sky130_fd_sc_hd__nor2_1 _26417_ (.A(_04245_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__nand2_1 _26418_ (.A(_04237_),
    .B(_04231_),
    .Y(_04248_));
 sky130_fd_sc_hd__or2_1 _26419_ (.A(_04247_),
    .B(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__nand2_1 _26420_ (.A(_04248_),
    .B(_04247_),
    .Y(_04250_));
 sky130_fd_sc_hd__a2bb2o_1 _26421_ (.A1_N(_01837_),
    .A2_N(_04149_),
    .B1(_04150_),
    .B2(_01832_),
    .X(_04251_));
 sky130_fd_sc_hd__nor2_1 _26422_ (.A(_01831_),
    .B(_04190_),
    .Y(_04252_));
 sky130_fd_sc_hd__a311o_1 _26423_ (.A1(_04249_),
    .A2(_04147_),
    .A3(_04250_),
    .B1(_04251_),
    .C1(_04252_),
    .X(_01838_));
 sky130_vsdinv _26424_ (.A(net34),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _26425_ (.A(_04223_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21a_1 _26426_ (.A1(_04225_),
    .A2(_01842_),
    .B1(_04227_),
    .X(_01843_));
 sky130_fd_sc_hd__nand2_1 _26427_ (.A(\count_instr[42] ),
    .B(_04167_),
    .Y(_04253_));
 sky130_fd_sc_hd__o221a_1 _26428_ (.A1(_19105_),
    .A2(_04180_),
    .B1(_04193_),
    .B2(_19416_),
    .C1(_04253_),
    .X(_01847_));
 sky130_fd_sc_hd__clkbuf_2 _26429_ (.A(_18713_),
    .X(_04254_));
 sky130_fd_sc_hd__a22o_1 _26430_ (.A1(\irq_mask[10] ),
    .A2(_04254_),
    .B1(_04243_),
    .B2(\timer[10] ),
    .X(_04255_));
 sky130_fd_sc_hd__a21oi_1 _26431_ (.A1(\cpuregs_rs1[10] ),
    .A2(_04141_),
    .B1(_04255_),
    .Y(_01849_));
 sky130_fd_sc_hd__buf_4 _26432_ (.A(_19316_),
    .X(_04256_));
 sky130_fd_sc_hd__o22ai_4 _26433_ (.A1(_01844_),
    .A2(_04120_),
    .B1(_04256_),
    .B2(_01850_),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_4 _26434_ (.A(_20722_),
    .B(_20645_),
    .Y(_04258_));
 sky130_vsdinv _26435_ (.A(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__and3_1 _26436_ (.A(_04247_),
    .B(_04231_),
    .C(_04230_),
    .X(_04260_));
 sky130_fd_sc_hd__o21ai_2 _26437_ (.A1(_04234_),
    .A2(_04235_),
    .B1(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__o21ba_1 _26438_ (.A1(_04231_),
    .A2(_04245_),
    .B1_N(_04246_),
    .X(_04262_));
 sky130_fd_sc_hd__nor2_2 _26439_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .Y(_04263_));
 sky130_fd_sc_hd__a21oi_4 _26440_ (.A1(_04261_),
    .A2(_04262_),
    .B1(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__or2_1 _26441_ (.A(_04263_),
    .B(_04258_),
    .X(_04265_));
 sky130_fd_sc_hd__a31o_1 _26442_ (.A1(_04261_),
    .A2(_04262_),
    .A3(_04265_),
    .B1(_18767_),
    .X(_04266_));
 sky130_fd_sc_hd__a21oi_2 _26443_ (.A1(_04259_),
    .A2(_04264_),
    .B1(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a211o_1 _26444_ (.A1(_20388_),
    .A2(_01845_),
    .B1(_04257_),
    .C1(_04267_),
    .X(_01851_));
 sky130_vsdinv _26445_ (.A(net35),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _26446_ (.A(_04223_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o21a_1 _26447_ (.A1(_04225_),
    .A2(_01855_),
    .B1(_04227_),
    .X(_01856_));
 sky130_fd_sc_hd__nand2_1 _26448_ (.A(\count_instr[11] ),
    .B(_20010_),
    .Y(_04268_));
 sky130_fd_sc_hd__o221a_1 _26449_ (.A1(_19160_),
    .A2(_04106_),
    .B1(_04193_),
    .B2(_19417_),
    .C1(_04268_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_2 _26450_ (.A(_04128_),
    .X(_04269_));
 sky130_fd_sc_hd__a22o_1 _26451_ (.A1(\irq_mask[11] ),
    .A2(_04254_),
    .B1(_04243_),
    .B2(\timer[11] ),
    .X(_04270_));
 sky130_fd_sc_hd__a21oi_1 _26452_ (.A1(\cpuregs_rs1[11] ),
    .A2(_04269_),
    .B1(_04270_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _26453_ (.A(_20732_),
    .B(_20646_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand2_2 _26454_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_1 _26455_ (.A(_04271_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__nor2_1 _26456_ (.A(_04258_),
    .B(_04264_),
    .Y(_04274_));
 sky130_fd_sc_hd__or2_1 _26457_ (.A(_04273_),
    .B(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__nand2_1 _26458_ (.A(_04274_),
    .B(_04273_),
    .Y(_04276_));
 sky130_fd_sc_hd__a2bb2o_1 _26459_ (.A1_N(_01863_),
    .A2_N(_04149_),
    .B1(_04150_),
    .B2(_01858_),
    .X(_04277_));
 sky130_fd_sc_hd__nor2_2 _26460_ (.A(_01857_),
    .B(_04190_),
    .Y(_04278_));
 sky130_fd_sc_hd__a311o_1 _26461_ (.A1(_04275_),
    .A2(_04147_),
    .A3(_04276_),
    .B1(_04277_),
    .C1(_04278_),
    .X(_01864_));
 sky130_vsdinv _26462_ (.A(net528),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _26463_ (.A(_04223_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__o21a_1 _26464_ (.A1(_04225_),
    .A2(_01868_),
    .B1(_04227_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_1 _26465_ (.A(_20012_),
    .B(\count_cycle[44] ),
    .Y(_04279_));
 sky130_fd_sc_hd__o221a_1 _26466_ (.A1(_19143_),
    .A2(_04106_),
    .B1(_19100_),
    .B2(_04108_),
    .C1(_04279_),
    .X(_01873_));
 sky130_fd_sc_hd__a22o_1 _26467_ (.A1(\irq_mask[12] ),
    .A2(_04254_),
    .B1(_04243_),
    .B2(\timer[12] ),
    .X(_04280_));
 sky130_fd_sc_hd__a21oi_1 _26468_ (.A1(\cpuregs_rs1[12] ),
    .A2(_04269_),
    .B1(_04280_),
    .Y(_01875_));
 sky130_fd_sc_hd__nor2_2 _26469_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .Y(_04281_));
 sky130_fd_sc_hd__nor2_2 _26470_ (.A(_20740_),
    .B(_20647_),
    .Y(_04282_));
 sky130_fd_sc_hd__nor2_1 _26471_ (.A(_04281_),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__o21ai_2 _26472_ (.A1(_04258_),
    .A2(_04264_),
    .B1(_04271_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_1 _26473_ (.A(_04284_),
    .B(_04272_),
    .Y(_04285_));
 sky130_fd_sc_hd__or2_1 _26474_ (.A(_04283_),
    .B(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__buf_2 _26475_ (.A(_18697_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_1 _26476_ (.A(_04285_),
    .B(_04283_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2_1 _26477_ (.A(_04122_),
    .B(_01871_),
    .Y(_04289_));
 sky130_fd_sc_hd__o221ai_4 _26478_ (.A1(_01870_),
    .A2(_04120_),
    .B1(_01876_),
    .B2(_04256_),
    .C1(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__a31o_1 _26479_ (.A1(_04286_),
    .A2(_04287_),
    .A3(_04288_),
    .B1(_04290_),
    .X(_01877_));
 sky130_vsdinv _26480_ (.A(net37),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _26481_ (.A(_04223_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21a_1 _26482_ (.A1(_04225_),
    .A2(_01881_),
    .B1(_04227_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_2 _26483_ (.A(_04105_),
    .X(_04291_));
 sky130_fd_sc_hd__nand2_1 _26484_ (.A(\count_instr[13] ),
    .B(_20010_),
    .Y(_04292_));
 sky130_fd_sc_hd__o221a_1 _26485_ (.A1(_19142_),
    .A2(_04291_),
    .B1(_04193_),
    .B2(_19458_),
    .C1(_04292_),
    .X(_01886_));
 sky130_fd_sc_hd__a22o_1 _26486_ (.A1(\irq_mask[13] ),
    .A2(_04254_),
    .B1(_04243_),
    .B2(\timer[13] ),
    .X(_04293_));
 sky130_fd_sc_hd__a21oi_1 _26487_ (.A1(\cpuregs_rs1[13] ),
    .A2(_04269_),
    .B1(_04293_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_1 _26488_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_04294_));
 sky130_fd_sc_hd__nor2_1 _26489_ (.A(_20746_),
    .B(_20648_),
    .Y(_04295_));
 sky130_fd_sc_hd__or2_1 _26490_ (.A(_04294_),
    .B(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__a21oi_2 _26491_ (.A1(_04284_),
    .A2(_04272_),
    .B1(_04281_),
    .Y(_04297_));
 sky130_fd_sc_hd__nor2_1 _26492_ (.A(_04282_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__or2_1 _26493_ (.A(_04296_),
    .B(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__nand2_1 _26494_ (.A(_04298_),
    .B(_04296_),
    .Y(_04300_));
 sky130_fd_sc_hd__a2bb2o_1 _26495_ (.A1_N(_01889_),
    .A2_N(_04149_),
    .B1(_04150_),
    .B2(_01884_),
    .X(_04301_));
 sky130_fd_sc_hd__nor2_2 _26496_ (.A(_01883_),
    .B(_04190_),
    .Y(_04302_));
 sky130_fd_sc_hd__a311o_1 _26497_ (.A1(_04299_),
    .A2(_04147_),
    .A3(_04300_),
    .B1(_04301_),
    .C1(_04302_),
    .X(_01890_));
 sky130_vsdinv _26498_ (.A(net38),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_1 _26499_ (.A(_04104_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21a_1 _26500_ (.A1(_04224_),
    .A2(_01894_),
    .B1(_04226_),
    .X(_01895_));
 sky130_vsdinv _26501_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_fd_sc_hd__nand2_1 _26502_ (.A(\count_instr[46] ),
    .B(_04167_),
    .Y(_04303_));
 sky130_fd_sc_hd__o221a_1 _26503_ (.A1(_19098_),
    .A2(_04180_),
    .B1(_04109_),
    .B2(_19459_),
    .C1(_04303_),
    .X(_01899_));
 sky130_fd_sc_hd__nand2_1 _26504_ (.A(\cpuregs_rs1[14] ),
    .B(_04129_),
    .Y(_04304_));
 sky130_fd_sc_hd__o221a_1 _26505_ (.A1(_18650_),
    .A2(_04114_),
    .B1(_04126_),
    .B2(_20574_),
    .C1(_04304_),
    .X(_01901_));
 sky130_fd_sc_hd__nor2_2 _26506_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .Y(_04305_));
 sky130_fd_sc_hd__nor2_4 _26507_ (.A(_20754_),
    .B(_20649_),
    .Y(_04306_));
 sky130_fd_sc_hd__or2_1 _26508_ (.A(_04305_),
    .B(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__o21bai_2 _26509_ (.A1(_04282_),
    .A2(_04297_),
    .B1_N(_04294_),
    .Y(_04308_));
 sky130_vsdinv _26510_ (.A(_04295_),
    .Y(_04309_));
 sky130_fd_sc_hd__and2_1 _26511_ (.A(_04308_),
    .B(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__or2_1 _26512_ (.A(_04307_),
    .B(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__nand2_1 _26513_ (.A(_04310_),
    .B(_04307_),
    .Y(_04312_));
 sky130_fd_sc_hd__o22a_1 _26514_ (.A1(_01896_),
    .A2(_04176_),
    .B1(_04239_),
    .B2(_01902_),
    .X(_04313_));
 sky130_fd_sc_hd__a21bo_1 _26515_ (.A1(_04204_),
    .A2(_01897_),
    .B1_N(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__a31o_1 _26516_ (.A1(_04311_),
    .A2(_04287_),
    .A3(_04312_),
    .B1(_04314_),
    .X(_01903_));
 sky130_vsdinv _26517_ (.A(net527),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _26518_ (.A(_04104_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o21a_4 _26519_ (.A1(_04224_),
    .A2(_01907_),
    .B1(_04226_),
    .X(_01908_));
 sky130_fd_sc_hd__nand2_1 _26520_ (.A(\count_instr[15] ),
    .B(_20010_),
    .Y(_04315_));
 sky130_fd_sc_hd__o221a_2 _26521_ (.A1(_19140_),
    .A2(_04291_),
    .B1(_04109_),
    .B2(_19457_),
    .C1(_04315_),
    .X(_01912_));
 sky130_fd_sc_hd__clkbuf_2 _26522_ (.A(_18714_),
    .X(_04316_));
 sky130_vsdinv _26523_ (.A(\timer[15] ),
    .Y(_04317_));
 sky130_fd_sc_hd__clkbuf_2 _26524_ (.A(_04128_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _26525_ (.A(\cpuregs_rs1[15] ),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__o221a_1 _26526_ (.A1(_18648_),
    .A2(_04316_),
    .B1(_04126_),
    .B2(_04317_),
    .C1(_04319_),
    .X(_01914_));
 sky130_fd_sc_hd__nor2_1 _26527_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .Y(_04320_));
 sky130_fd_sc_hd__nor2_2 _26528_ (.A(_20759_),
    .B(_20650_),
    .Y(_04321_));
 sky130_fd_sc_hd__or2_2 _26529_ (.A(_04320_),
    .B(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__a21oi_4 _26530_ (.A1(_04308_),
    .A2(_04309_),
    .B1(_04305_),
    .Y(_04323_));
 sky130_fd_sc_hd__nor2_4 _26531_ (.A(_04306_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__nor2_4 _26532_ (.A(_04322_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__a21o_1 _26533_ (.A1(_04324_),
    .A2(_04322_),
    .B1(_20539_),
    .X(_04326_));
 sky130_fd_sc_hd__o2bb2a_1 _26534_ (.A1_N(_04122_),
    .A2_N(_01910_),
    .B1(_01915_),
    .B2(_04205_),
    .X(_04327_));
 sky130_fd_sc_hd__o221ai_2 _26535_ (.A1(_20541_),
    .A2(_01909_),
    .B1(_04325_),
    .B2(_04326_),
    .C1(_04327_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_1 _26536_ (.A(net450),
    .B(net40),
    .Y(_01917_));
 sky130_fd_sc_hd__clkbuf_2 _26537_ (.A(instr_rdcycleh),
    .X(_04328_));
 sky130_fd_sc_hd__nand2_1 _26538_ (.A(_04328_),
    .B(\count_cycle[48] ),
    .Y(_04329_));
 sky130_fd_sc_hd__o221a_2 _26539_ (.A1(_19139_),
    .A2(_04291_),
    .B1(_19097_),
    .B2(_04108_),
    .C1(_04329_),
    .X(_01921_));
 sky130_fd_sc_hd__a22o_1 _26540_ (.A1(\irq_mask[16] ),
    .A2(_04254_),
    .B1(_04243_),
    .B2(\timer[16] ),
    .X(_04330_));
 sky130_fd_sc_hd__a21oi_1 _26541_ (.A1(\cpuregs_rs1[16] ),
    .A2(_04269_),
    .B1(_04330_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _26542_ (.A(_20767_),
    .B(_20652_),
    .Y(_04331_));
 sky130_vsdinv _26543_ (.A(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_1 _26544_ (.A(_20767_),
    .B(_20652_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand2_1 _26545_ (.A(_04332_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__nor2_1 _26546_ (.A(_04321_),
    .B(_04325_),
    .Y(_04335_));
 sky130_fd_sc_hd__nor2_1 _26547_ (.A(_04334_),
    .B(_04335_),
    .Y(_04336_));
 sky130_vsdinv _26548_ (.A(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _26549_ (.A(_04335_),
    .B(_04334_),
    .Y(_04338_));
 sky130_fd_sc_hd__a2bb2o_1 _26550_ (.A1_N(_01924_),
    .A2_N(_04205_),
    .B1(_20387_),
    .B2(_01919_),
    .X(_04339_));
 sky130_fd_sc_hd__nor2_4 _26551_ (.A(_01918_),
    .B(_04190_),
    .Y(_04340_));
 sky130_fd_sc_hd__a311o_1 _26552_ (.A1(_04337_),
    .A2(_04147_),
    .A3(_04338_),
    .B1(_04339_),
    .C1(_04340_),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_1 _26553_ (.A(net450),
    .B(net41),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _26554_ (.A(\count_instr[49] ),
    .B(_20005_),
    .Y(_04341_));
 sky130_fd_sc_hd__o221a_2 _26555_ (.A1(_19273_),
    .A2(_04180_),
    .B1(_04109_),
    .B2(_19496_),
    .C1(_04341_),
    .X(_01930_));
 sky130_fd_sc_hd__clkbuf_2 _26556_ (.A(_19974_),
    .X(_04342_));
 sky130_fd_sc_hd__a22o_1 _26557_ (.A1(\irq_mask[17] ),
    .A2(_04254_),
    .B1(_04342_),
    .B2(\timer[17] ),
    .X(_04343_));
 sky130_fd_sc_hd__a21oi_1 _26558_ (.A1(\cpuregs_rs1[17] ),
    .A2(_04269_),
    .B1(_04343_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_2 _26559_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_04344_));
 sky130_fd_sc_hd__nor2_2 _26560_ (.A(_20772_),
    .B(_20653_),
    .Y(_04345_));
 sky130_fd_sc_hd__nor2_1 _26561_ (.A(_04344_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand2_1 _26562_ (.A(_04337_),
    .B(_04332_),
    .Y(_04347_));
 sky130_fd_sc_hd__or2_1 _26563_ (.A(_04346_),
    .B(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__nand2_1 _26564_ (.A(_04347_),
    .B(_04346_),
    .Y(_04349_));
 sky130_fd_sc_hd__a2bb2o_1 _26565_ (.A1_N(_01933_),
    .A2_N(_04205_),
    .B1(_20387_),
    .B2(_01928_),
    .X(_04350_));
 sky130_fd_sc_hd__nor2_4 _26566_ (.A(_01927_),
    .B(_04190_),
    .Y(_04351_));
 sky130_fd_sc_hd__a311o_1 _26567_ (.A1(_04348_),
    .A2(_04349_),
    .A3(_04116_),
    .B1(_04350_),
    .C1(_04351_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_1 _26568_ (.A(net450),
    .B(net42),
    .Y(_01935_));
 sky130_fd_sc_hd__clkbuf_2 _26569_ (.A(instr_rdcycleh),
    .X(_04352_));
 sky130_fd_sc_hd__a22o_1 _26570_ (.A1(\count_instr[18] ),
    .A2(_20009_),
    .B1(_04352_),
    .B2(\count_cycle[50] ),
    .X(_04353_));
 sky130_fd_sc_hd__a21oi_4 _26571_ (.A1(\count_instr[50] ),
    .A2(_20006_),
    .B1(_04353_),
    .Y(_01939_));
 sky130_fd_sc_hd__clkbuf_2 _26572_ (.A(_18712_),
    .X(_04354_));
 sky130_fd_sc_hd__nand2_1 _26573_ (.A(\cpuregs_rs1[18] ),
    .B(_04318_),
    .Y(_04355_));
 sky130_fd_sc_hd__o221a_1 _26574_ (.A1(_18608_),
    .A2(_04316_),
    .B1(_04354_),
    .B2(_20579_),
    .C1(_04355_),
    .X(_01941_));
 sky130_fd_sc_hd__nor2_2 _26575_ (.A(\reg_pc[18] ),
    .B(_20654_),
    .Y(_04356_));
 sky130_fd_sc_hd__nor2_2 _26576_ (.A(\decoded_imm[18] ),
    .B(_20779_),
    .Y(_04357_));
 sky130_fd_sc_hd__o21ba_1 _26577_ (.A1(_04344_),
    .A2(_04332_),
    .B1_N(_04345_),
    .X(_04358_));
 sky130_vsdinv _26578_ (.A(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__o21bai_2 _26579_ (.A1(_04306_),
    .A2(_04323_),
    .B1_N(_04320_),
    .Y(_04360_));
 sky130_vsdinv _26580_ (.A(_04321_),
    .Y(_04361_));
 sky130_fd_sc_hd__or3_4 _26581_ (.A(_04344_),
    .B(_04345_),
    .C(_04334_),
    .X(_04362_));
 sky130_fd_sc_hd__a21oi_4 _26582_ (.A1(_04360_),
    .A2(_04361_),
    .B1(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__or4_4 _26583_ (.A(_04356_),
    .B(_04357_),
    .C(_04359_),
    .D(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__o22ai_4 _26584_ (.A1(_04356_),
    .A2(_04357_),
    .B1(_04359_),
    .B2(_04363_),
    .Y(_04365_));
 sky130_fd_sc_hd__o22ai_1 _26585_ (.A1(_01936_),
    .A2(_04119_),
    .B1(_04205_),
    .B2(_01942_),
    .Y(_04366_));
 sky130_fd_sc_hd__a21o_1 _26586_ (.A1(_04136_),
    .A2(_01937_),
    .B1(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__a31o_1 _26587_ (.A1(_04364_),
    .A2(_04287_),
    .A3(_04365_),
    .B1(_04367_),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_1 _26588_ (.A(net450),
    .B(net526),
    .Y(_01944_));
 sky130_vsdinv _26589_ (.A(\count_cycle[19] ),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _26590_ (.A(_04328_),
    .B(\count_cycle[51] ),
    .Y(_04368_));
 sky130_fd_sc_hd__o221a_1 _26591_ (.A1(_19148_),
    .A2(_04291_),
    .B1(_19122_),
    .B2(_04108_),
    .C1(_04368_),
    .X(_01948_));
 sky130_fd_sc_hd__nand2_1 _26592_ (.A(\cpuregs_rs1[19] ),
    .B(_04318_),
    .Y(_04369_));
 sky130_fd_sc_hd__o221a_1 _26593_ (.A1(_18606_),
    .A2(_04316_),
    .B1(_04354_),
    .B2(_20578_),
    .C1(_04369_),
    .X(_01950_));
 sky130_fd_sc_hd__nand2_1 _26594_ (.A(_20788_),
    .B(\decoded_imm[19] ),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_2 _26595_ (.A(_20655_),
    .B(\reg_pc[19] ),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_2 _26596_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .Y(_04372_));
 sky130_fd_sc_hd__a22oi_4 _26597_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04365_),
    .B2(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__and4_1 _26598_ (.A(_04365_),
    .B(_04372_),
    .C(_04370_),
    .D(_04371_),
    .X(_04374_));
 sky130_fd_sc_hd__o22a_2 _26599_ (.A1(_01945_),
    .A2(_18960_),
    .B1(_04149_),
    .B2(_01951_),
    .X(_04375_));
 sky130_fd_sc_hd__nand2_1 _26600_ (.A(_20388_),
    .B(_01946_),
    .Y(_04376_));
 sky130_fd_sc_hd__o311ai_1 _26601_ (.A1(_20540_),
    .A2(_04373_),
    .A3(_04374_),
    .B1(_04375_),
    .C1(_04376_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand2_1 _26602_ (.A(net450),
    .B(net524),
    .Y(_01953_));
 sky130_fd_sc_hd__clkbuf_2 _26603_ (.A(_04107_),
    .X(_04377_));
 sky130_fd_sc_hd__nand2_1 _26604_ (.A(_04328_),
    .B(\count_cycle[52] ),
    .Y(_04378_));
 sky130_fd_sc_hd__o221a_1 _26605_ (.A1(_19147_),
    .A2(_04291_),
    .B1(_19121_),
    .B2(_04377_),
    .C1(_04378_),
    .X(_01957_));
 sky130_fd_sc_hd__clkbuf_2 _26606_ (.A(_18713_),
    .X(_04379_));
 sky130_fd_sc_hd__a22o_1 _26607_ (.A1(\irq_mask[20] ),
    .A2(_04379_),
    .B1(_04342_),
    .B2(\timer[20] ),
    .X(_04380_));
 sky130_fd_sc_hd__a21oi_4 _26608_ (.A1(\cpuregs_rs1[20] ),
    .A2(_04269_),
    .B1(_04380_),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_1 _26609_ (.A(_20794_),
    .B(_20656_),
    .Y(_04381_));
 sky130_vsdinv _26610_ (.A(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _26611_ (.A(_20794_),
    .B(_20656_),
    .Y(_04383_));
 sky130_fd_sc_hd__nand2_1 _26612_ (.A(_04382_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__nor2_2 _26613_ (.A(_20788_),
    .B(_20655_),
    .Y(_04385_));
 sky130_fd_sc_hd__or2_1 _26614_ (.A(_04385_),
    .B(_04373_),
    .X(_04386_));
 sky130_vsdinv _26615_ (.A(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__or2_1 _26616_ (.A(_04384_),
    .B(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_1 _26617_ (.A(_04387_),
    .B(_04384_),
    .Y(_04389_));
 sky130_fd_sc_hd__o22a_1 _26618_ (.A1(_01954_),
    .A2(_04176_),
    .B1(_04239_),
    .B2(_01960_),
    .X(_04390_));
 sky130_fd_sc_hd__a21bo_2 _26619_ (.A1(_04204_),
    .A2(_01955_),
    .B1_N(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__a31o_1 _26620_ (.A1(_04388_),
    .A2(_04287_),
    .A3(_04389_),
    .B1(_04391_),
    .X(_01961_));
 sky130_fd_sc_hd__clkbuf_2 _26621_ (.A(_04093_),
    .X(_04392_));
 sky130_fd_sc_hd__nand2_1 _26622_ (.A(_04392_),
    .B(net46),
    .Y(_01962_));
 sky130_fd_sc_hd__nand2_1 _26623_ (.A(\count_instr[21] ),
    .B(_20010_),
    .Y(_04393_));
 sky130_fd_sc_hd__o221a_1 _26624_ (.A1(_19197_),
    .A2(_04291_),
    .B1(_04109_),
    .B2(_19408_),
    .C1(_04393_),
    .X(_01966_));
 sky130_fd_sc_hd__buf_4 _26625_ (.A(_04128_),
    .X(_04394_));
 sky130_fd_sc_hd__a22o_1 _26626_ (.A1(\irq_mask[21] ),
    .A2(_04379_),
    .B1(_04342_),
    .B2(\timer[21] ),
    .X(_04395_));
 sky130_fd_sc_hd__a21oi_4 _26627_ (.A1(\cpuregs_rs1[21] ),
    .A2(_04394_),
    .B1(_04395_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_2 _26628_ (.A(_20802_),
    .B(_20657_),
    .Y(_04396_));
 sky130_vsdinv _26629_ (.A(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _26630_ (.A(_20802_),
    .B(_20657_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _26631_ (.A(_04397_),
    .B(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__o22ai_4 _26632_ (.A1(\reg_pc[20] ),
    .A2(\decoded_imm[20] ),
    .B1(_04385_),
    .B2(_04373_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _26633_ (.A(_04400_),
    .B(_04382_),
    .Y(_04401_));
 sky130_vsdinv _26634_ (.A(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__or2_1 _26635_ (.A(_04399_),
    .B(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__nand2_1 _26636_ (.A(_04402_),
    .B(_04399_),
    .Y(_04404_));
 sky130_fd_sc_hd__o22a_1 _26637_ (.A1(_01963_),
    .A2(_04176_),
    .B1(_04239_),
    .B2(_01969_),
    .X(_04405_));
 sky130_fd_sc_hd__a21bo_2 _26638_ (.A1(_04204_),
    .A2(_01964_),
    .B1_N(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__a31o_1 _26639_ (.A1(_04403_),
    .A2(_04287_),
    .A3(_04404_),
    .B1(_04406_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _26640_ (.A(_04392_),
    .B(net47),
    .Y(_01971_));
 sky130_fd_sc_hd__a22o_1 _26641_ (.A1(\count_instr[54] ),
    .A2(_20005_),
    .B1(\count_instr[22] ),
    .B2(_20009_),
    .X(_04407_));
 sky130_fd_sc_hd__a21oi_1 _26642_ (.A1(_20012_),
    .A2(\count_cycle[54] ),
    .B1(_04407_),
    .Y(_01975_));
 sky130_fd_sc_hd__a22o_1 _26643_ (.A1(\irq_mask[22] ),
    .A2(_04379_),
    .B1(_04342_),
    .B2(\timer[22] ),
    .X(_04408_));
 sky130_fd_sc_hd__a21oi_4 _26644_ (.A1(\cpuregs_rs1[22] ),
    .A2(_04394_),
    .B1(_04408_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _26645_ (.A(_20807_),
    .B(_20659_),
    .Y(_04409_));
 sky130_vsdinv _26646_ (.A(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nor2_1 _26647_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .Y(_04411_));
 sky130_vsdinv _26648_ (.A(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2_1 _26649_ (.A(_04410_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__a22oi_4 _26650_ (.A1(_20802_),
    .A2(_20657_),
    .B1(_04400_),
    .B2(_04382_),
    .Y(_04414_));
 sky130_vsdinv _26651_ (.A(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_1 _26652_ (.A(_04415_),
    .B(_04397_),
    .Y(_04416_));
 sky130_vsdinv _26653_ (.A(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__or2_1 _26654_ (.A(_04413_),
    .B(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__nand2_1 _26655_ (.A(_04417_),
    .B(_04413_),
    .Y(_04419_));
 sky130_fd_sc_hd__o22a_1 _26656_ (.A1(_01972_),
    .A2(_04176_),
    .B1(_04239_),
    .B2(_01978_),
    .X(_04420_));
 sky130_fd_sc_hd__a21bo_2 _26657_ (.A1(_04204_),
    .A2(_01973_),
    .B1_N(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__a31o_1 _26658_ (.A1(_04418_),
    .A2(_04287_),
    .A3(_04419_),
    .B1(_04421_),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_1 _26659_ (.A(_04392_),
    .B(net48),
    .Y(_01980_));
 sky130_fd_sc_hd__clkbuf_2 _26660_ (.A(_04105_),
    .X(_04422_));
 sky130_fd_sc_hd__nand2_1 _26661_ (.A(_04328_),
    .B(\count_cycle[55] ),
    .Y(_04423_));
 sky130_fd_sc_hd__o221a_1 _26662_ (.A1(_19192_),
    .A2(_04422_),
    .B1(_19259_),
    .B2(_04377_),
    .C1(_04423_),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_1 _26663_ (.A1(\irq_mask[23] ),
    .A2(_04379_),
    .B1(_04342_),
    .B2(\timer[23] ),
    .X(_04424_));
 sky130_fd_sc_hd__a21oi_4 _26664_ (.A1(\cpuregs_rs1[23] ),
    .A2(_04394_),
    .B1(_04424_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _26665_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_4 _26666_ (.A(_20815_),
    .B(_20660_),
    .Y(_04426_));
 sky130_fd_sc_hd__or2_1 _26667_ (.A(_04425_),
    .B(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__o22ai_4 _26668_ (.A1(\reg_pc[22] ),
    .A2(\decoded_imm[22] ),
    .B1(_04396_),
    .B2(_04414_),
    .Y(_04428_));
 sky130_fd_sc_hd__and2_1 _26669_ (.A(_04428_),
    .B(_04410_),
    .X(_04429_));
 sky130_fd_sc_hd__or2_1 _26670_ (.A(_04427_),
    .B(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__nand2_1 _26671_ (.A(_04429_),
    .B(_04427_),
    .Y(_04431_));
 sky130_fd_sc_hd__o22a_1 _26672_ (.A1(_01981_),
    .A2(_18722_),
    .B1(_04239_),
    .B2(_01987_),
    .X(_04432_));
 sky130_fd_sc_hd__a21bo_2 _26673_ (.A1(_04204_),
    .A2(_01982_),
    .B1_N(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__a31o_1 _26674_ (.A1(_04430_),
    .A2(_04116_),
    .A3(_04431_),
    .B1(_04433_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _26675_ (.A(_04392_),
    .B(net49),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _26676_ (.A(_04328_),
    .B(\count_cycle[56] ),
    .Y(_04434_));
 sky130_fd_sc_hd__o221a_1 _26677_ (.A1(_19186_),
    .A2(_04422_),
    .B1(_19265_),
    .B2(_04377_),
    .C1(_04434_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_1 _26678_ (.A(\cpuregs_rs1[24] ),
    .B(_04318_),
    .Y(_04435_));
 sky130_fd_sc_hd__o221a_1 _26679_ (.A1(_18614_),
    .A2(_04316_),
    .B1(_04354_),
    .B2(_20626_),
    .C1(_04435_),
    .X(_01995_));
 sky130_fd_sc_hd__nand2_1 _26680_ (.A(_20821_),
    .B(_20661_),
    .Y(_04436_));
 sky130_fd_sc_hd__nand2_2 _26681_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _26682_ (.A(_04436_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__a22oi_4 _26683_ (.A1(_20815_),
    .A2(_20660_),
    .B1(_04428_),
    .B2(_04410_),
    .Y(_04439_));
 sky130_fd_sc_hd__nor2_1 _26684_ (.A(_04426_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__or2_1 _26685_ (.A(_04438_),
    .B(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__nand2_1 _26686_ (.A(_04440_),
    .B(_04438_),
    .Y(_04442_));
 sky130_fd_sc_hd__o22ai_1 _26687_ (.A1(_01990_),
    .A2(_04119_),
    .B1(_19316_),
    .B2(_01996_),
    .Y(_04443_));
 sky130_fd_sc_hd__a21o_2 _26688_ (.A1(_04136_),
    .A2(_01991_),
    .B1(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__a31o_1 _26689_ (.A1(_04441_),
    .A2(_04116_),
    .A3(_04442_),
    .B1(_04444_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _26690_ (.A(_04392_),
    .B(net50),
    .Y(_01998_));
 sky130_vsdinv _26691_ (.A(\count_cycle[25] ),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2_1 _26692_ (.A(_04328_),
    .B(\count_cycle[57] ),
    .Y(_04445_));
 sky130_fd_sc_hd__o221a_1 _26693_ (.A1(_19183_),
    .A2(_04422_),
    .B1(_19096_),
    .B2(_04377_),
    .C1(_04445_),
    .X(_02002_));
 sky130_fd_sc_hd__a22o_1 _26694_ (.A1(\irq_mask[25] ),
    .A2(_04379_),
    .B1(_04342_),
    .B2(\timer[25] ),
    .X(_04446_));
 sky130_fd_sc_hd__a21oi_4 _26695_ (.A1(\cpuregs_rs1[25] ),
    .A2(_04394_),
    .B1(_04446_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _26696_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_04447_));
 sky130_fd_sc_hd__nor2_1 _26697_ (.A(_20827_),
    .B(_20662_),
    .Y(_04448_));
 sky130_fd_sc_hd__or2_1 _26698_ (.A(_04447_),
    .B(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__a21o_1 _26699_ (.A1(_04441_),
    .A2(_04437_),
    .B1(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__a31oi_1 _26700_ (.A1(_04441_),
    .A2(_04437_),
    .A3(_04449_),
    .B1(_20539_),
    .Y(_04451_));
 sky130_fd_sc_hd__o22ai_4 _26701_ (.A1(_01999_),
    .A2(_04120_),
    .B1(_04256_),
    .B2(_02005_),
    .Y(_04452_));
 sky130_fd_sc_hd__a221o_1 _26702_ (.A1(_20388_),
    .A2(_02000_),
    .B1(_04450_),
    .B2(_04451_),
    .C1(_04452_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2_1 _26703_ (.A(_04392_),
    .B(net51),
    .Y(_02007_));
 sky130_fd_sc_hd__a22o_1 _26704_ (.A1(\count_instr[58] ),
    .A2(_20005_),
    .B1(\count_instr[26] ),
    .B2(_20009_),
    .X(_04453_));
 sky130_fd_sc_hd__a21oi_2 _26705_ (.A1(_20012_),
    .A2(\count_cycle[58] ),
    .B1(_04453_),
    .Y(_02011_));
 sky130_fd_sc_hd__a22o_1 _26706_ (.A1(\irq_mask[26] ),
    .A2(_04379_),
    .B1(_19974_),
    .B2(\timer[26] ),
    .X(_04454_));
 sky130_fd_sc_hd__a21oi_1 _26707_ (.A1(\cpuregs_rs1[26] ),
    .A2(_04394_),
    .B1(_04454_),
    .Y(_02013_));
 sky130_fd_sc_hd__o2bb2a_1 _26708_ (.A1_N(_04122_),
    .A2_N(_02009_),
    .B1(_02014_),
    .B2(_04205_),
    .X(_04455_));
 sky130_fd_sc_hd__or2_1 _26709_ (.A(_04438_),
    .B(_04449_),
    .X(_04456_));
 sky130_fd_sc_hd__o21bai_4 _26710_ (.A1(_04426_),
    .A2(_04439_),
    .B1_N(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__o21ba_1 _26711_ (.A1(_04437_),
    .A2(_04447_),
    .B1_N(_04448_),
    .X(_04458_));
 sky130_fd_sc_hd__nor2_1 _26712_ (.A(_20833_),
    .B(_20663_),
    .Y(_04459_));
 sky130_vsdinv _26713_ (.A(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _26714_ (.A(_20833_),
    .B(_20663_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_1 _26715_ (.A(_04460_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__a21oi_1 _26716_ (.A1(_04457_),
    .A2(_04458_),
    .B1(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__and3_1 _26717_ (.A(_04457_),
    .B(_04458_),
    .C(_04462_),
    .X(_04464_));
 sky130_fd_sc_hd__or3_4 _26718_ (.A(_20539_),
    .B(_04463_),
    .C(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__o211ai_2 _26719_ (.A1(_20541_),
    .A2(_02008_),
    .B1(_04455_),
    .C1(_04465_),
    .Y(_02015_));
 sky130_fd_sc_hd__clkbuf_2 _26720_ (.A(_04093_),
    .X(_04466_));
 sky130_fd_sc_hd__nand2_1 _26721_ (.A(_04466_),
    .B(net52),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_1 _26722_ (.A(_04352_),
    .B(\count_cycle[59] ),
    .Y(_04467_));
 sky130_fd_sc_hd__o221a_1 _26723_ (.A1(_19155_),
    .A2(_04422_),
    .B1(_19127_),
    .B2(_04377_),
    .C1(_04467_),
    .X(_02020_));
 sky130_fd_sc_hd__a22o_1 _26724_ (.A1(\irq_mask[27] ),
    .A2(_18713_),
    .B1(_19974_),
    .B2(\timer[27] ),
    .X(_04468_));
 sky130_fd_sc_hd__a21oi_2 _26725_ (.A1(\cpuregs_rs1[27] ),
    .A2(_04394_),
    .B1(_04468_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_2 _26726_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_04469_));
 sky130_fd_sc_hd__nor2_2 _26727_ (.A(_20843_),
    .B(_20664_),
    .Y(_04470_));
 sky130_fd_sc_hd__nor2_1 _26728_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__or2_1 _26729_ (.A(_04459_),
    .B(_04463_),
    .X(_04472_));
 sky130_fd_sc_hd__or2_1 _26730_ (.A(_04471_),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__nand2_1 _26731_ (.A(_04472_),
    .B(_04471_),
    .Y(_04474_));
 sky130_fd_sc_hd__o2bb2a_1 _26732_ (.A1_N(_20387_),
    .A2_N(_02018_),
    .B1(_02023_),
    .B2(_19335_),
    .X(_04475_));
 sky130_fd_sc_hd__o21ai_2 _26733_ (.A1(_04120_),
    .A2(_02017_),
    .B1(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__a31o_1 _26734_ (.A1(_04473_),
    .A2(_04116_),
    .A3(_04474_),
    .B1(_04476_),
    .X(_02024_));
 sky130_fd_sc_hd__nand2_1 _26735_ (.A(_04466_),
    .B(net53),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _26736_ (.A(_04352_),
    .B(_19472_),
    .Y(_04477_));
 sky130_fd_sc_hd__o221a_1 _26737_ (.A1(_19154_),
    .A2(_04422_),
    .B1(_19131_),
    .B2(_04377_),
    .C1(_04477_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _26738_ (.A(\cpuregs_rs1[28] ),
    .B(_04318_),
    .Y(_04478_));
 sky130_fd_sc_hd__o221a_1 _26739_ (.A1(_18638_),
    .A2(_04316_),
    .B1(_04354_),
    .B2(_20633_),
    .C1(_04478_),
    .X(_02031_));
 sky130_fd_sc_hd__nor2_1 _26740_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_04479_));
 sky130_fd_sc_hd__nor2_1 _26741_ (.A(_20848_),
    .B(_20665_),
    .Y(_04480_));
 sky130_fd_sc_hd__nor2_1 _26742_ (.A(_04479_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__o21ba_1 _26743_ (.A1(_04469_),
    .A2(_04460_),
    .B1_N(_04470_),
    .X(_04482_));
 sky130_vsdinv _26744_ (.A(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__or3_4 _26745_ (.A(_04469_),
    .B(_04470_),
    .C(_04462_),
    .X(_04484_));
 sky130_fd_sc_hd__a21oi_4 _26746_ (.A1(_04457_),
    .A2(_04458_),
    .B1(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__or2_1 _26747_ (.A(_04483_),
    .B(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__or2_1 _26748_ (.A(_04481_),
    .B(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__nand2_1 _26749_ (.A(_04486_),
    .B(_04481_),
    .Y(_04488_));
 sky130_fd_sc_hd__o22ai_4 _26750_ (.A1(_02026_),
    .A2(_18960_),
    .B1(_19317_),
    .B2(_02032_),
    .Y(_04489_));
 sky130_fd_sc_hd__and2_1 _26751_ (.A(_04122_),
    .B(_02027_),
    .X(_04490_));
 sky130_fd_sc_hd__a311o_1 _26752_ (.A1(_04487_),
    .A2(_18697_),
    .A3(_04488_),
    .B1(_04489_),
    .C1(_04490_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_1 _26753_ (.A(_04466_),
    .B(net54),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _26754_ (.A(_04352_),
    .B(\count_cycle[61] ),
    .Y(_04491_));
 sky130_fd_sc_hd__o221a_1 _26755_ (.A1(_19169_),
    .A2(_04422_),
    .B1(_19130_),
    .B2(_04111_),
    .C1(_04491_),
    .X(_02038_));
 sky130_fd_sc_hd__a22o_1 _26756_ (.A1(\irq_mask[29] ),
    .A2(_18713_),
    .B1(_19974_),
    .B2(\timer[29] ),
    .X(_04492_));
 sky130_fd_sc_hd__a21oi_1 _26757_ (.A1(\cpuregs_rs1[29] ),
    .A2(_04129_),
    .B1(_04492_),
    .Y(_02040_));
 sky130_vsdinv _26758_ (.A(_02036_),
    .Y(_04493_));
 sky130_fd_sc_hd__o22ai_4 _26759_ (.A1(\reg_pc[28] ),
    .A2(\decoded_imm[28] ),
    .B1(_04483_),
    .B2(_04485_),
    .Y(_04494_));
 sky130_vsdinv _26760_ (.A(_04480_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_2 _26761_ (.A(_20857_),
    .B(_20666_),
    .Y(_04496_));
 sky130_vsdinv _26762_ (.A(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__nand2_1 _26763_ (.A(_20857_),
    .B(_20666_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _26764_ (.A(_04497_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__a21oi_1 _26765_ (.A1(_04494_),
    .A2(_04495_),
    .B1(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__a31o_1 _26766_ (.A1(_04494_),
    .A2(_04495_),
    .A3(_04499_),
    .B1(_20539_),
    .X(_04501_));
 sky130_fd_sc_hd__o22a_1 _26767_ (.A1(_02035_),
    .A2(_18960_),
    .B1(_19324_),
    .B2(_02041_),
    .X(_04502_));
 sky130_fd_sc_hd__o221ai_1 _26768_ (.A1(_18743_),
    .A2(_04493_),
    .B1(_04500_),
    .B2(_04501_),
    .C1(_04502_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _26769_ (.A(_04466_),
    .B(net523),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _26770_ (.A(_04352_),
    .B(\count_cycle[62] ),
    .Y(_04503_));
 sky130_fd_sc_hd__o221a_1 _26771_ (.A1(_19168_),
    .A2(_04105_),
    .B1(_19129_),
    .B2(_04111_),
    .C1(_04503_),
    .X(_02047_));
 sky130_vsdinv _26772_ (.A(\timer[30] ),
    .Y(_04504_));
 sky130_fd_sc_hd__nand2_1 _26773_ (.A(\cpuregs_rs1[30] ),
    .B(_04318_),
    .Y(_04505_));
 sky130_fd_sc_hd__o221a_1 _26774_ (.A1(_18642_),
    .A2(_04316_),
    .B1(_04354_),
    .B2(_04504_),
    .C1(_04505_),
    .X(_02049_));
 sky130_fd_sc_hd__a22oi_4 _26775_ (.A1(_20857_),
    .A2(_20666_),
    .B1(_04494_),
    .B2(_04495_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_2 _26776_ (.A(\reg_pc[30] ),
    .B(_20667_),
    .Y(_04507_));
 sky130_fd_sc_hd__nor2_2 _26777_ (.A(\decoded_imm[30] ),
    .B(_20864_),
    .Y(_04508_));
 sky130_fd_sc_hd__nor2_1 _26778_ (.A(_04507_),
    .B(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand3b_1 _26779_ (.A_N(_04506_),
    .B(_04497_),
    .C(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__o22ai_4 _26780_ (.A1(_04507_),
    .A2(_04508_),
    .B1(_04496_),
    .B2(_04506_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_2 _26781_ (.A(_02050_),
    .B(_04256_),
    .Y(_04512_));
 sky130_fd_sc_hd__a2bb2o_1 _26782_ (.A1_N(_02044_),
    .A2_N(_18960_),
    .B1(_04150_),
    .B2(_02045_),
    .X(_04513_));
 sky130_fd_sc_hd__a311o_1 _26783_ (.A1(_04510_),
    .A2(_04511_),
    .A3(_04116_),
    .B1(_04512_),
    .C1(_04513_),
    .X(_02051_));
 sky130_fd_sc_hd__nand2_1 _26784_ (.A(_04466_),
    .B(net57),
    .Y(_02052_));
 sky130_fd_sc_hd__a22o_1 _26785_ (.A1(\count_instr[31] ),
    .A2(_20009_),
    .B1(_04352_),
    .B2(\count_cycle[63] ),
    .X(_04514_));
 sky130_fd_sc_hd__a21oi_2 _26786_ (.A1(\count_instr[63] ),
    .A2(_20006_),
    .B1(_04514_),
    .Y(_02056_));
 sky130_vsdinv _26787_ (.A(\timer[31] ),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _26788_ (.A(\cpuregs_rs1[31] ),
    .B(_04128_),
    .Y(_04516_));
 sky130_fd_sc_hd__o221a_1 _26789_ (.A1(_18640_),
    .A2(_18714_),
    .B1(_04354_),
    .B2(_04515_),
    .C1(_04516_),
    .X(_02058_));
 sky130_fd_sc_hd__nand2_1 _26790_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .Y(_04517_));
 sky130_fd_sc_hd__xnor2_1 _26791_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_1 _26792_ (.A1(_04511_),
    .A2(_04517_),
    .B1(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__nand3_1 _26793_ (.A(_04511_),
    .B(_04517_),
    .C(_04518_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _26794_ (.A(_04520_),
    .B(_18697_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_1 _26795_ (.A(_04122_),
    .B(_02054_),
    .Y(_04522_));
 sky130_fd_sc_hd__o221ai_4 _26796_ (.A1(_02053_),
    .A2(_04120_),
    .B1(_02059_),
    .B2(_04256_),
    .C1(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__o21bai_1 _26797_ (.A1(_04519_),
    .A2(_04521_),
    .B1_N(_04523_),
    .Y(_02060_));
 sky130_fd_sc_hd__or2_1 _26798_ (.A(\decoded_rd[4] ),
    .B(_00308_),
    .X(_02061_));
 sky130_vsdinv _26799_ (.A(_20367_),
    .Y(_02062_));
 sky130_fd_sc_hd__o21ai_1 _26800_ (.A1(_02064_),
    .A2(_20540_),
    .B1(_04256_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor3_2 _26801_ (.A(_18661_),
    .B(_02410_),
    .C(_00308_),
    .Y(_02066_));
 sky130_fd_sc_hd__and3_1 _26802_ (.A(_18959_),
    .B(_20540_),
    .C(_20541_),
    .X(_02067_));
 sky130_fd_sc_hd__nand2_1 _26803_ (.A(_18699_),
    .B(_00343_),
    .Y(_04524_));
 sky130_fd_sc_hd__a211o_1 _26804_ (.A1(_04524_),
    .A2(_20390_),
    .B1(_18704_),
    .C1(_18544_),
    .X(_02068_));
 sky130_fd_sc_hd__nor2_4 _26805_ (.A(latched_branch),
    .B(_18746_),
    .Y(_04525_));
 sky130_fd_sc_hd__clkbuf_2 _26806_ (.A(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_4 _26807_ (.A(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__nor2_4 _26808_ (.A(_04527_),
    .B(_19596_),
    .Y(_02069_));
 sky130_fd_sc_hd__clkbuf_2 _26809_ (.A(_18754_),
    .X(_04528_));
 sky130_fd_sc_hd__nor2_1 _26810_ (.A(_18749_),
    .B(_20669_),
    .Y(_04529_));
 sky130_fd_sc_hd__a221o_1 _26811_ (.A1(_18597_),
    .A2(_04528_),
    .B1(_04527_),
    .B2(_02070_),
    .C1(_04529_),
    .X(_02071_));
 sky130_fd_sc_hd__and2_1 _26812_ (.A(_18761_),
    .B(\reg_next_pc[1] ),
    .X(_04530_));
 sky130_fd_sc_hd__a221o_1 _26813_ (.A1(_18599_),
    .A2(_04528_),
    .B1(_04527_),
    .B2(_01465_),
    .C1(_04530_),
    .X(_02072_));
 sky130_fd_sc_hd__clkbuf_4 _26814_ (.A(_04526_),
    .X(_04531_));
 sky130_fd_sc_hd__and3_1 _26815_ (.A(_18595_),
    .B(_18759_),
    .C(\irq_pending[2] ),
    .X(_04532_));
 sky130_fd_sc_hd__a221o_1 _26816_ (.A1(_20878_),
    .A2(\reg_next_pc[2] ),
    .B1(_00293_),
    .B2(_04531_),
    .C1(_04532_),
    .X(_02074_));
 sky130_fd_sc_hd__nor2_1 _26817_ (.A(\reg_pc[3] ),
    .B(\reg_pc[2] ),
    .Y(_04533_));
 sky130_fd_sc_hd__nor2_2 _26818_ (.A(_19087_),
    .B(_02073_),
    .Y(_04534_));
 sky130_fd_sc_hd__nor2_1 _26819_ (.A(_04533_),
    .B(_04534_),
    .Y(_02075_));
 sky130_fd_sc_hd__buf_2 _26820_ (.A(_04526_),
    .X(_04535_));
 sky130_fd_sc_hd__and3_1 _26821_ (.A(_18600_),
    .B(_18759_),
    .C(\irq_pending[3] ),
    .X(_04536_));
 sky130_fd_sc_hd__a221o_1 _26822_ (.A1(_20878_),
    .A2(\reg_next_pc[3] ),
    .B1(_01468_),
    .B2(_04535_),
    .C1(_04536_),
    .X(_02076_));
 sky130_fd_sc_hd__nor2_1 _26823_ (.A(\reg_pc[4] ),
    .B(_04534_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _26824_ (.A(_04534_),
    .B(\reg_pc[4] ),
    .Y(_04538_));
 sky130_vsdinv _26825_ (.A(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_2 _26826_ (.A(_04537_),
    .B(_04539_),
    .Y(_02077_));
 sky130_fd_sc_hd__and3_1 _26827_ (.A(_18634_),
    .B(_18759_),
    .C(\irq_pending[4] ),
    .X(_04540_));
 sky130_fd_sc_hd__a221o_1 _26828_ (.A1(_20878_),
    .A2(\reg_next_pc[4] ),
    .B1(_01472_),
    .B2(_04535_),
    .C1(_04540_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_2 _26829_ (.A(_20688_),
    .B(_04538_),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_1 _26830_ (.A(\reg_pc[5] ),
    .B(_04539_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_2 _26831_ (.A(_04541_),
    .B(_04542_),
    .Y(_02079_));
 sky130_fd_sc_hd__and3_1 _26832_ (.A(_18633_),
    .B(_18759_),
    .C(\irq_pending[5] ),
    .X(_04543_));
 sky130_fd_sc_hd__a221o_1 _26833_ (.A1(_20878_),
    .A2(\reg_next_pc[5] ),
    .B1(_01476_),
    .B2(_04535_),
    .C1(_04543_),
    .X(_02080_));
 sky130_fd_sc_hd__nor2_1 _26834_ (.A(\reg_pc[6] ),
    .B(_04541_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _26835_ (.A(_04541_),
    .B(\reg_pc[6] ),
    .Y(_04545_));
 sky130_vsdinv _26836_ (.A(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__nor2_1 _26837_ (.A(_04544_),
    .B(_04546_),
    .Y(_02081_));
 sky130_fd_sc_hd__buf_2 _26838_ (.A(\irq_state[0] ),
    .X(_04547_));
 sky130_fd_sc_hd__and2_1 _26839_ (.A(_04547_),
    .B(\reg_next_pc[6] ),
    .X(_04548_));
 sky130_fd_sc_hd__a221o_2 _26840_ (.A1(_18632_),
    .A2(_04528_),
    .B1(_04527_),
    .B2(_01479_),
    .C1(_04548_),
    .X(_02082_));
 sky130_fd_sc_hd__nor2_2 _26841_ (.A(_20701_),
    .B(_04545_),
    .Y(_04549_));
 sky130_fd_sc_hd__nor2_1 _26842_ (.A(\reg_pc[7] ),
    .B(_04546_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _26843_ (.A(_04549_),
    .B(_04550_),
    .Y(_02083_));
 sky130_fd_sc_hd__and2_1 _26844_ (.A(_04547_),
    .B(\reg_next_pc[7] ),
    .X(_04551_));
 sky130_fd_sc_hd__a221o_2 _26845_ (.A1(_18631_),
    .A2(_04528_),
    .B1(_04527_),
    .B2(_01482_),
    .C1(_04551_),
    .X(_02084_));
 sky130_fd_sc_hd__or2_1 _26846_ (.A(\reg_pc[8] ),
    .B(_04549_),
    .X(_04552_));
 sky130_fd_sc_hd__nand2_1 _26847_ (.A(_04549_),
    .B(\reg_pc[8] ),
    .Y(_04553_));
 sky130_fd_sc_hd__and2_1 _26848_ (.A(_04552_),
    .B(_04553_),
    .X(_02085_));
 sky130_fd_sc_hd__and3_1 _26849_ (.A(_18628_),
    .B(_18759_),
    .C(\irq_pending[8] ),
    .X(_04554_));
 sky130_fd_sc_hd__a221o_1 _26850_ (.A1(_20878_),
    .A2(\reg_next_pc[8] ),
    .B1(_01485_),
    .B2(_04535_),
    .C1(_04554_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_2 _26851_ (.A(_20716_),
    .B(_04553_),
    .Y(_04555_));
 sky130_fd_sc_hd__and2_1 _26852_ (.A(_04553_),
    .B(_20716_),
    .X(_04556_));
 sky130_fd_sc_hd__nor2_1 _26853_ (.A(_04555_),
    .B(_04556_),
    .Y(_02087_));
 sky130_fd_sc_hd__clkbuf_4 _26854_ (.A(_18761_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_2 _26855_ (.A(\irq_state[1] ),
    .X(_04558_));
 sky130_fd_sc_hd__and3_1 _26856_ (.A(_18627_),
    .B(_04558_),
    .C(\irq_pending[9] ),
    .X(_04559_));
 sky130_fd_sc_hd__a221o_1 _26857_ (.A1(_04557_),
    .A2(\reg_next_pc[9] ),
    .B1(_01488_),
    .B2(_04535_),
    .C1(_04559_),
    .X(_02088_));
 sky130_fd_sc_hd__nor2_1 _26858_ (.A(\reg_pc[10] ),
    .B(_04555_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _26859_ (.A(_04555_),
    .B(\reg_pc[10] ),
    .Y(_04561_));
 sky130_vsdinv _26860_ (.A(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__nor2_1 _26861_ (.A(_04560_),
    .B(_04562_),
    .Y(_02089_));
 sky130_fd_sc_hd__and2_1 _26862_ (.A(_04547_),
    .B(\reg_next_pc[10] ),
    .X(_04563_));
 sky130_fd_sc_hd__a221o_2 _26863_ (.A1(_18626_),
    .A2(_04528_),
    .B1(_04527_),
    .B2(_01491_),
    .C1(_04563_),
    .X(_02090_));
 sky130_fd_sc_hd__nor2_2 _26864_ (.A(_20732_),
    .B(_04561_),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _26865_ (.A(\reg_pc[11] ),
    .B(_04562_),
    .Y(_04565_));
 sky130_fd_sc_hd__nor2_1 _26866_ (.A(_04564_),
    .B(_04565_),
    .Y(_02091_));
 sky130_fd_sc_hd__and2_1 _26867_ (.A(_04547_),
    .B(\reg_next_pc[11] ),
    .X(_04566_));
 sky130_fd_sc_hd__a221o_2 _26868_ (.A1(_18625_),
    .A2(_04528_),
    .B1(_04531_),
    .B2(_01494_),
    .C1(_04566_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _26869_ (.A(\reg_pc[12] ),
    .B(_04564_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand2_1 _26870_ (.A(_04564_),
    .B(\reg_pc[12] ),
    .Y(_04568_));
 sky130_vsdinv _26871_ (.A(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_1 _26872_ (.A(_04567_),
    .B(_04569_),
    .Y(_02093_));
 sky130_fd_sc_hd__and3_1 _26873_ (.A(_18646_),
    .B(_04558_),
    .C(\irq_pending[12] ),
    .X(_04570_));
 sky130_fd_sc_hd__a221o_1 _26874_ (.A1(_04557_),
    .A2(\reg_next_pc[12] ),
    .B1(_01497_),
    .B2(_04535_),
    .C1(_04570_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_2 _26875_ (.A(_20746_),
    .B(_04568_),
    .Y(_04571_));
 sky130_fd_sc_hd__nor2_1 _26876_ (.A(\reg_pc[13] ),
    .B(_04569_),
    .Y(_04572_));
 sky130_fd_sc_hd__nor2_1 _26877_ (.A(_04571_),
    .B(_04572_),
    .Y(_02095_));
 sky130_fd_sc_hd__clkbuf_4 _26878_ (.A(_04525_),
    .X(_04573_));
 sky130_fd_sc_hd__and3_1 _26879_ (.A(_18645_),
    .B(_04558_),
    .C(\irq_pending[13] ),
    .X(_04574_));
 sky130_fd_sc_hd__a221o_1 _26880_ (.A1(_04557_),
    .A2(\reg_next_pc[13] ),
    .B1(_01500_),
    .B2(_04573_),
    .C1(_04574_),
    .X(_02096_));
 sky130_fd_sc_hd__nor2_1 _26881_ (.A(\reg_pc[14] ),
    .B(_04571_),
    .Y(_04575_));
 sky130_fd_sc_hd__and2_1 _26882_ (.A(_04571_),
    .B(\reg_pc[14] ),
    .X(_04576_));
 sky130_fd_sc_hd__nor2_1 _26883_ (.A(_04575_),
    .B(_04576_),
    .Y(_02097_));
 sky130_fd_sc_hd__and3_1 _26884_ (.A(_18650_),
    .B(_04558_),
    .C(\irq_pending[14] ),
    .X(_04577_));
 sky130_fd_sc_hd__a221o_1 _26885_ (.A1(_04557_),
    .A2(\reg_next_pc[14] ),
    .B1(_01503_),
    .B2(_04573_),
    .C1(_04577_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_1 _26886_ (.A(\reg_pc[15] ),
    .B(_04576_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _26887_ (.A(_04576_),
    .B(\reg_pc[15] ),
    .Y(_04579_));
 sky130_vsdinv _26888_ (.A(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__nor2_1 _26889_ (.A(_04578_),
    .B(_04580_),
    .Y(_02099_));
 sky130_fd_sc_hd__and3_2 _26890_ (.A(_18648_),
    .B(_04558_),
    .C(\irq_pending[15] ),
    .X(_04581_));
 sky130_fd_sc_hd__a221o_1 _26891_ (.A1(_04557_),
    .A2(\reg_next_pc[15] ),
    .B1(_01506_),
    .B2(_04573_),
    .C1(_04581_),
    .X(_02100_));
 sky130_fd_sc_hd__nor2_2 _26892_ (.A(_20767_),
    .B(_04579_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _26893_ (.A(\reg_pc[16] ),
    .B(_04580_),
    .Y(_04583_));
 sky130_fd_sc_hd__nor2_1 _26894_ (.A(_04582_),
    .B(_04583_),
    .Y(_02101_));
 sky130_fd_sc_hd__and2_1 _26895_ (.A(_04547_),
    .B(\reg_next_pc[16] ),
    .X(_04584_));
 sky130_fd_sc_hd__a221o_1 _26896_ (.A1(_18605_),
    .A2(_18754_),
    .B1(_04531_),
    .B2(_01509_),
    .C1(_04584_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_1 _26897_ (.A(\reg_pc[17] ),
    .B(_04582_),
    .Y(_04585_));
 sky130_fd_sc_hd__and2_1 _26898_ (.A(_04582_),
    .B(\reg_pc[17] ),
    .X(_04586_));
 sky130_fd_sc_hd__nor2_1 _26899_ (.A(_04585_),
    .B(_04586_),
    .Y(_02103_));
 sky130_fd_sc_hd__and3_1 _26900_ (.A(_18603_),
    .B(_04558_),
    .C(\irq_pending[17] ),
    .X(_04587_));
 sky130_fd_sc_hd__a221o_1 _26901_ (.A1(_04557_),
    .A2(\reg_next_pc[17] ),
    .B1(_01512_),
    .B2(_04573_),
    .C1(_04587_),
    .X(_02104_));
 sky130_fd_sc_hd__or2_1 _26902_ (.A(\reg_pc[18] ),
    .B(_04586_),
    .X(_04588_));
 sky130_fd_sc_hd__nand2_1 _26903_ (.A(_04586_),
    .B(\reg_pc[18] ),
    .Y(_04589_));
 sky130_fd_sc_hd__and2_1 _26904_ (.A(_04588_),
    .B(_04589_),
    .X(_02105_));
 sky130_fd_sc_hd__buf_2 _26905_ (.A(_18761_),
    .X(_04590_));
 sky130_fd_sc_hd__buf_1 _26906_ (.A(\irq_state[1] ),
    .X(_04591_));
 sky130_fd_sc_hd__and3_1 _26907_ (.A(_18608_),
    .B(_04591_),
    .C(\irq_pending[18] ),
    .X(_04592_));
 sky130_fd_sc_hd__a221o_1 _26908_ (.A1(_04590_),
    .A2(\reg_next_pc[18] ),
    .B1(_01515_),
    .B2(_04573_),
    .C1(_04592_),
    .X(_02106_));
 sky130_fd_sc_hd__nor2_1 _26909_ (.A(_20788_),
    .B(_04589_),
    .Y(_04593_));
 sky130_fd_sc_hd__and2_1 _26910_ (.A(_04589_),
    .B(_20788_),
    .X(_04594_));
 sky130_fd_sc_hd__nor2_1 _26911_ (.A(_04593_),
    .B(_04594_),
    .Y(_02107_));
 sky130_fd_sc_hd__and3_1 _26912_ (.A(_18606_),
    .B(_04591_),
    .C(\irq_pending[19] ),
    .X(_04595_));
 sky130_fd_sc_hd__a221o_1 _26913_ (.A1(_04590_),
    .A2(\reg_next_pc[19] ),
    .B1(_01518_),
    .B2(_04573_),
    .C1(_04595_),
    .X(_02108_));
 sky130_fd_sc_hd__nor2_1 _26914_ (.A(\reg_pc[20] ),
    .B(_04593_),
    .Y(_04596_));
 sky130_fd_sc_hd__and2_1 _26915_ (.A(_04593_),
    .B(\reg_pc[20] ),
    .X(_04597_));
 sky130_fd_sc_hd__nor2_1 _26916_ (.A(_04596_),
    .B(_04597_),
    .Y(_02109_));
 sky130_fd_sc_hd__buf_2 _26917_ (.A(_04525_),
    .X(_04598_));
 sky130_fd_sc_hd__and3_1 _26918_ (.A(_18621_),
    .B(_04591_),
    .C(\irq_pending[20] ),
    .X(_04599_));
 sky130_fd_sc_hd__a221o_1 _26919_ (.A1(_04590_),
    .A2(\reg_next_pc[20] ),
    .B1(_01521_),
    .B2(_04598_),
    .C1(_04599_),
    .X(_02110_));
 sky130_fd_sc_hd__or2_1 _26920_ (.A(\reg_pc[21] ),
    .B(_04597_),
    .X(_04600_));
 sky130_fd_sc_hd__nand2_1 _26921_ (.A(_04597_),
    .B(\reg_pc[21] ),
    .Y(_04601_));
 sky130_fd_sc_hd__and2_1 _26922_ (.A(_04600_),
    .B(_04601_),
    .X(_02111_));
 sky130_fd_sc_hd__and3_1 _26923_ (.A(_18620_),
    .B(_04591_),
    .C(\irq_pending[21] ),
    .X(_04602_));
 sky130_fd_sc_hd__a221o_1 _26924_ (.A1(_04590_),
    .A2(\reg_next_pc[21] ),
    .B1(_01524_),
    .B2(_04598_),
    .C1(_04602_),
    .X(_02112_));
 sky130_fd_sc_hd__nor2_2 _26925_ (.A(_20807_),
    .B(_04601_),
    .Y(_04603_));
 sky130_fd_sc_hd__and2_1 _26926_ (.A(_04601_),
    .B(_20807_),
    .X(_04604_));
 sky130_fd_sc_hd__nor2_1 _26927_ (.A(_04603_),
    .B(_04604_),
    .Y(_02113_));
 sky130_fd_sc_hd__and2_1 _26928_ (.A(_04547_),
    .B(\reg_next_pc[22] ),
    .X(_04605_));
 sky130_fd_sc_hd__a221o_1 _26929_ (.A1(_18619_),
    .A2(_18754_),
    .B1(_04531_),
    .B2(_01527_),
    .C1(_04605_),
    .X(_02114_));
 sky130_fd_sc_hd__or2_1 _26930_ (.A(\reg_pc[23] ),
    .B(_04603_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2_1 _26931_ (.A(_04603_),
    .B(\reg_pc[23] ),
    .Y(_04607_));
 sky130_fd_sc_hd__and2_1 _26932_ (.A(_04606_),
    .B(_04607_),
    .X(_02115_));
 sky130_fd_sc_hd__and3_1 _26933_ (.A(_18617_),
    .B(_04591_),
    .C(\irq_pending[23] ),
    .X(_04608_));
 sky130_fd_sc_hd__a221o_1 _26934_ (.A1(_04590_),
    .A2(\reg_next_pc[23] ),
    .B1(_01530_),
    .B2(_04598_),
    .C1(_04608_),
    .X(_02116_));
 sky130_fd_sc_hd__nor2_2 _26935_ (.A(_20821_),
    .B(_04607_),
    .Y(_04609_));
 sky130_fd_sc_hd__and2_1 _26936_ (.A(_04607_),
    .B(_20821_),
    .X(_04610_));
 sky130_fd_sc_hd__nor2_1 _26937_ (.A(_04609_),
    .B(_04610_),
    .Y(_02117_));
 sky130_fd_sc_hd__and3_1 _26938_ (.A(_18614_),
    .B(_04591_),
    .C(\irq_pending[24] ),
    .X(_04611_));
 sky130_fd_sc_hd__a221o_1 _26939_ (.A1(_04590_),
    .A2(\reg_next_pc[24] ),
    .B1(_01533_),
    .B2(_04598_),
    .C1(_04611_),
    .X(_02118_));
 sky130_fd_sc_hd__nor2_1 _26940_ (.A(\reg_pc[25] ),
    .B(_04609_),
    .Y(_04612_));
 sky130_fd_sc_hd__nand2_1 _26941_ (.A(_04609_),
    .B(\reg_pc[25] ),
    .Y(_04613_));
 sky130_vsdinv _26942_ (.A(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_1 _26943_ (.A(_04612_),
    .B(_04614_),
    .Y(_02119_));
 sky130_fd_sc_hd__and3_1 _26944_ (.A(_18613_),
    .B(_18753_),
    .C(\irq_pending[25] ),
    .X(_04615_));
 sky130_fd_sc_hd__a221o_1 _26945_ (.A1(_18762_),
    .A2(\reg_next_pc[25] ),
    .B1(_01536_),
    .B2(_04598_),
    .C1(_04615_),
    .X(_02120_));
 sky130_fd_sc_hd__nor2_2 _26946_ (.A(_20833_),
    .B(_04613_),
    .Y(_04616_));
 sky130_fd_sc_hd__nor2_1 _26947_ (.A(\reg_pc[26] ),
    .B(_04614_),
    .Y(_04617_));
 sky130_fd_sc_hd__nor2_1 _26948_ (.A(_04616_),
    .B(_04617_),
    .Y(_02121_));
 sky130_fd_sc_hd__and2_1 _26949_ (.A(_18748_),
    .B(\reg_next_pc[26] ),
    .X(_04618_));
 sky130_fd_sc_hd__a221o_1 _26950_ (.A1(_18612_),
    .A2(_18754_),
    .B1(_04531_),
    .B2(_01539_),
    .C1(_04618_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_1 _26951_ (.A(\reg_pc[27] ),
    .B(_04616_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _26952_ (.A(_04616_),
    .B(\reg_pc[27] ),
    .Y(_04620_));
 sky130_vsdinv _26953_ (.A(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__nor2_1 _26954_ (.A(_04619_),
    .B(_04621_),
    .Y(_02123_));
 sky130_fd_sc_hd__and2_1 _26955_ (.A(_18748_),
    .B(\reg_next_pc[27] ),
    .X(_04622_));
 sky130_fd_sc_hd__a221o_1 _26956_ (.A1(_18611_),
    .A2(_18754_),
    .B1(_04531_),
    .B2(_01542_),
    .C1(_04622_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_2 _26957_ (.A(_20848_),
    .B(_04620_),
    .Y(_04623_));
 sky130_fd_sc_hd__nor2_1 _26958_ (.A(\reg_pc[28] ),
    .B(_04621_),
    .Y(_04624_));
 sky130_fd_sc_hd__nor2_1 _26959_ (.A(_04623_),
    .B(_04624_),
    .Y(_02125_));
 sky130_fd_sc_hd__and3_1 _26960_ (.A(_18638_),
    .B(_18753_),
    .C(\irq_pending[28] ),
    .X(_04625_));
 sky130_fd_sc_hd__a221o_1 _26961_ (.A1(_18762_),
    .A2(\reg_next_pc[28] ),
    .B1(_01545_),
    .B2(_04598_),
    .C1(_04625_),
    .X(_02126_));
 sky130_fd_sc_hd__nor2_1 _26962_ (.A(\reg_pc[29] ),
    .B(_04623_),
    .Y(_04626_));
 sky130_fd_sc_hd__and2_1 _26963_ (.A(_04623_),
    .B(\reg_pc[29] ),
    .X(_04627_));
 sky130_fd_sc_hd__nor2_1 _26964_ (.A(_04626_),
    .B(_04627_),
    .Y(_02127_));
 sky130_fd_sc_hd__and3_1 _26965_ (.A(_18637_),
    .B(_18753_),
    .C(\irq_pending[29] ),
    .X(_04628_));
 sky130_fd_sc_hd__a221o_1 _26966_ (.A1(_18762_),
    .A2(\reg_next_pc[29] ),
    .B1(_01548_),
    .B2(_04526_),
    .C1(_04628_),
    .X(_02128_));
 sky130_fd_sc_hd__or2_1 _26967_ (.A(\reg_pc[30] ),
    .B(_04627_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _26968_ (.A(_04627_),
    .B(\reg_pc[30] ),
    .Y(_04630_));
 sky130_fd_sc_hd__and2_1 _26969_ (.A(_04629_),
    .B(_04630_),
    .X(_02129_));
 sky130_fd_sc_hd__and3_1 _26970_ (.A(_18642_),
    .B(_18753_),
    .C(\irq_pending[30] ),
    .X(_04631_));
 sky130_fd_sc_hd__a221o_1 _26971_ (.A1(_18762_),
    .A2(\reg_next_pc[30] ),
    .B1(_01551_),
    .B2(_04526_),
    .C1(_04631_),
    .X(_02130_));
 sky130_fd_sc_hd__xor2_1 _26972_ (.A(_20870_),
    .B(_04630_),
    .X(_02131_));
 sky130_fd_sc_hd__and3_1 _26973_ (.A(_18640_),
    .B(_18753_),
    .C(\irq_pending[31] ),
    .X(_04632_));
 sky130_fd_sc_hd__a221o_1 _26974_ (.A1(_18762_),
    .A2(\reg_next_pc[31] ),
    .B1(_01554_),
    .B2(_04526_),
    .C1(_04632_),
    .X(_02132_));
 sky130_fd_sc_hd__buf_2 _26975_ (.A(_18740_),
    .X(_04633_));
 sky130_vsdinv _26976_ (.A(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__nor2_8 _26977_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_04635_));
 sky130_fd_sc_hd__nor2_8 _26978_ (.A(instr_xor),
    .B(instr_xori),
    .Y(_04636_));
 sky130_fd_sc_hd__buf_2 _26979_ (.A(_04636_),
    .X(_04637_));
 sky130_vsdinv _26980_ (.A(is_compare),
    .Y(_04638_));
 sky130_fd_sc_hd__and3_1 _26981_ (.A(_04635_),
    .B(_04637_),
    .C(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__nor2_1 _26982_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04640_));
 sky130_vsdinv _26983_ (.A(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__nor2_8 _26984_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04642_));
 sky130_vsdinv _26985_ (.A(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__nor2_1 _26986_ (.A(_04641_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__and3_4 _26987_ (.A(_04634_),
    .B(_04639_),
    .C(_04644_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_2 _26988_ (.A(_18740_),
    .X(_04645_));
 sky130_fd_sc_hd__buf_2 _26989_ (.A(_04645_),
    .X(_04646_));
 sky130_vsdinv _26990_ (.A(_04636_),
    .Y(_04647_));
 sky130_fd_sc_hd__buf_2 _26991_ (.A(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__buf_2 _26992_ (.A(_04648_),
    .X(_04649_));
 sky130_vsdinv _26993_ (.A(_04635_),
    .Y(_04650_));
 sky130_fd_sc_hd__buf_2 _26994_ (.A(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__buf_2 _26995_ (.A(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__a21oi_1 _26996_ (.A1(_20392_),
    .A2(_20323_),
    .B1(_04642_),
    .Y(_04653_));
 sky130_vsdinv _26997_ (.A(_00343_),
    .Y(_04654_));
 sky130_fd_sc_hd__a32o_1 _26998_ (.A1(_04641_),
    .A2(_19677_),
    .A3(_20064_),
    .B1(_04654_),
    .B2(is_compare),
    .X(_04655_));
 sky130_fd_sc_hd__a211o_1 _26999_ (.A1(\alu_shl[0] ),
    .A2(_04652_),
    .B1(_04653_),
    .C1(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__a221o_1 _27000_ (.A1(\alu_shr[0] ),
    .A2(_04646_),
    .B1(_02591_),
    .B2(_04649_),
    .C1(_04656_),
    .X(_02134_));
 sky130_fd_sc_hd__buf_2 _27001_ (.A(_04650_),
    .X(_04657_));
 sky130_fd_sc_hd__buf_2 _27002_ (.A(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__buf_2 _27003_ (.A(_04643_),
    .X(_04659_));
 sky130_fd_sc_hd__buf_2 _27004_ (.A(_04659_),
    .X(_04660_));
 sky130_vsdinv _27005_ (.A(_04644_),
    .Y(_04661_));
 sky130_fd_sc_hd__buf_2 _27006_ (.A(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__o211a_1 _27007_ (.A1(_04660_),
    .A2(_20493_),
    .B1(_20495_),
    .C1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__nor2_1 _27008_ (.A(_04637_),
    .B(_20496_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21o_1 _27009_ (.A1(\alu_shr[1] ),
    .A2(_04633_),
    .B1(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__a211o_1 _27010_ (.A1(\alu_shl[1] ),
    .A2(_04658_),
    .B1(_04663_),
    .C1(_04665_),
    .X(_02135_));
 sky130_vsdinv _27011_ (.A(_20481_),
    .Y(_04666_));
 sky130_fd_sc_hd__buf_2 _27012_ (.A(_04660_),
    .X(_04667_));
 sky130_fd_sc_hd__buf_2 _27013_ (.A(_04641_),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_4 _27014_ (.A(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__buf_2 _27015_ (.A(_18740_),
    .X(_04670_));
 sky130_fd_sc_hd__a22o_1 _27016_ (.A1(_20484_),
    .A2(_04647_),
    .B1(_04670_),
    .B2(\alu_shr[2] ),
    .X(_04671_));
 sky130_fd_sc_hd__a21o_1 _27017_ (.A1(\alu_shl[2] ),
    .A2(_04658_),
    .B1(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__a221o_1 _27018_ (.A1(_04666_),
    .A2(_04667_),
    .B1(_20483_),
    .B2(_04669_),
    .C1(_04672_),
    .X(_02136_));
 sky130_vsdinv _27019_ (.A(_20477_),
    .Y(_04673_));
 sky130_fd_sc_hd__and2_1 _27020_ (.A(_04651_),
    .B(\alu_shl[3] ),
    .X(_04674_));
 sky130_fd_sc_hd__a221o_1 _27021_ (.A1(_20480_),
    .A2(_04647_),
    .B1(_04645_),
    .B2(\alu_shr[3] ),
    .C1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__a221o_1 _27022_ (.A1(_04673_),
    .A2(_04667_),
    .B1(_20479_),
    .B2(_04669_),
    .C1(_04675_),
    .X(_02137_));
 sky130_vsdinv _27023_ (.A(_20487_),
    .Y(_04676_));
 sky130_fd_sc_hd__nor2_1 _27024_ (.A(_04636_),
    .B(_20491_),
    .Y(_04677_));
 sky130_fd_sc_hd__a221o_1 _27025_ (.A1(\alu_shr[4] ),
    .A2(_04670_),
    .B1(\alu_shl[4] ),
    .B2(_04657_),
    .C1(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__a221o_1 _27026_ (.A1(_04676_),
    .A2(_04667_),
    .B1(_20489_),
    .B2(_04668_),
    .C1(_04678_),
    .X(_02138_));
 sky130_fd_sc_hd__or2_1 _27027_ (.A(_20470_),
    .B(_04659_),
    .X(_04679_));
 sky130_vsdinv _27028_ (.A(_20468_),
    .Y(_04680_));
 sky130_fd_sc_hd__a32o_1 _27029_ (.A1(_04662_),
    .A2(_04679_),
    .A3(_04680_),
    .B1(\alu_shl[5] ),
    .B2(_04652_),
    .X(_04681_));
 sky130_fd_sc_hd__a221o_1 _27030_ (.A1(\alu_shr[5] ),
    .A2(_04646_),
    .B1(_20471_),
    .B2(_04649_),
    .C1(_04681_),
    .X(_02139_));
 sky130_fd_sc_hd__or2_1 _27031_ (.A(_20473_),
    .B(_04659_),
    .X(_04682_));
 sky130_fd_sc_hd__a32o_1 _27032_ (.A1(_04662_),
    .A2(_20474_),
    .A3(_04682_),
    .B1(\alu_shl[6] ),
    .B2(_04652_),
    .X(_04683_));
 sky130_fd_sc_hd__a221o_1 _27033_ (.A1(\alu_shr[6] ),
    .A2(_04646_),
    .B1(_20476_),
    .B2(_04649_),
    .C1(_04683_),
    .X(_02140_));
 sky130_fd_sc_hd__inv_2 _27034_ (.A(net229),
    .Y(_02336_));
 sky130_fd_sc_hd__a21oi_1 _27035_ (.A1(_02336_),
    .A2(_20703_),
    .B1(_04642_),
    .Y(_04684_));
 sky130_fd_sc_hd__a21o_1 _27036_ (.A1(\alu_shl[7] ),
    .A2(_04652_),
    .B1(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__a2bb2o_1 _27037_ (.A1_N(_20497_),
    .A2_N(_04637_),
    .B1(\alu_shr[7] ),
    .B2(_04645_),
    .X(_04686_));
 sky130_fd_sc_hd__a311o_1 _27038_ (.A1(_19670_),
    .A2(_20057_),
    .A3(_04669_),
    .B1(_04685_),
    .C1(_04686_),
    .X(_02141_));
 sky130_vsdinv _27039_ (.A(_20459_),
    .Y(_04687_));
 sky130_fd_sc_hd__a22o_1 _27040_ (.A1(\alu_shl[8] ),
    .A2(_04657_),
    .B1(_04670_),
    .B2(\alu_shr[8] ),
    .X(_04688_));
 sky130_fd_sc_hd__a221o_1 _27041_ (.A1(_04687_),
    .A2(_04660_),
    .B1(_20462_),
    .B2(_04648_),
    .C1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__a21o_1 _27042_ (.A1(_20461_),
    .A2(_04669_),
    .B1(_04689_),
    .X(_02142_));
 sky130_fd_sc_hd__or2_1 _27043_ (.A(_20457_),
    .B(_04659_),
    .X(_04690_));
 sky130_vsdinv _27044_ (.A(_20455_),
    .Y(_04691_));
 sky130_fd_sc_hd__a32o_1 _27045_ (.A1(_04662_),
    .A2(_04690_),
    .A3(_04691_),
    .B1(\alu_shl[9] ),
    .B2(_04652_),
    .X(_04692_));
 sky130_fd_sc_hd__a221o_1 _27046_ (.A1(\alu_shr[9] ),
    .A2(_04646_),
    .B1(_20458_),
    .B2(_04649_),
    .C1(_04692_),
    .X(_02143_));
 sky130_fd_sc_hd__buf_2 _27047_ (.A(_04645_),
    .X(_04693_));
 sky130_fd_sc_hd__buf_2 _27048_ (.A(_04661_),
    .X(_04694_));
 sky130_fd_sc_hd__or2_1 _27049_ (.A(_20465_),
    .B(_04659_),
    .X(_04695_));
 sky130_vsdinv _27050_ (.A(_20463_),
    .Y(_04696_));
 sky130_fd_sc_hd__buf_2 _27051_ (.A(_04651_),
    .X(_04697_));
 sky130_fd_sc_hd__a32o_1 _27052_ (.A1(_04694_),
    .A2(_04695_),
    .A3(_04696_),
    .B1(\alu_shl[10] ),
    .B2(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__a221o_1 _27053_ (.A1(\alu_shr[10] ),
    .A2(_04693_),
    .B1(_20466_),
    .B2(_04649_),
    .C1(_04698_),
    .X(_02144_));
 sky130_vsdinv _27054_ (.A(_20451_),
    .Y(_04699_));
 sky130_fd_sc_hd__a22o_1 _27055_ (.A1(_20454_),
    .A2(_04647_),
    .B1(_04670_),
    .B2(\alu_shr[11] ),
    .X(_04700_));
 sky130_fd_sc_hd__a21o_1 _27056_ (.A1(\alu_shl[11] ),
    .A2(_04658_),
    .B1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__a221o_1 _27057_ (.A1(_04699_),
    .A2(_04667_),
    .B1(_20453_),
    .B2(_04668_),
    .C1(_04701_),
    .X(_02145_));
 sky130_vsdinv _27058_ (.A(_20435_),
    .Y(_04702_));
 sky130_fd_sc_hd__nor2_1 _27059_ (.A(_04636_),
    .B(_20439_),
    .Y(_04703_));
 sky130_fd_sc_hd__a221o_1 _27060_ (.A1(\alu_shl[12] ),
    .A2(_04657_),
    .B1(_04645_),
    .B2(\alu_shr[12] ),
    .C1(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__a221o_1 _27061_ (.A1(_04702_),
    .A2(_04667_),
    .B1(_20437_),
    .B2(_04668_),
    .C1(_04704_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_2 _27062_ (.A(_04643_),
    .X(_04705_));
 sky130_fd_sc_hd__or2_1 _27063_ (.A(_20432_),
    .B(_04705_),
    .X(_04706_));
 sky130_vsdinv _27064_ (.A(_20430_),
    .Y(_04707_));
 sky130_fd_sc_hd__a32o_1 _27065_ (.A1(_04694_),
    .A2(_04706_),
    .A3(_04707_),
    .B1(\alu_shl[13] ),
    .B2(_04697_),
    .X(_04708_));
 sky130_fd_sc_hd__a221o_1 _27066_ (.A1(\alu_shr[13] ),
    .A2(_04693_),
    .B1(_20433_),
    .B2(_04649_),
    .C1(_04708_),
    .X(_02147_));
 sky130_fd_sc_hd__buf_2 _27067_ (.A(_04648_),
    .X(_04709_));
 sky130_fd_sc_hd__or2_1 _27068_ (.A(_20442_),
    .B(_04705_),
    .X(_04710_));
 sky130_vsdinv _27069_ (.A(_20440_),
    .Y(_04711_));
 sky130_fd_sc_hd__a32o_1 _27070_ (.A1(_04694_),
    .A2(_04710_),
    .A3(_04711_),
    .B1(\alu_shl[14] ),
    .B2(_04697_),
    .X(_04712_));
 sky130_fd_sc_hd__a221o_1 _27071_ (.A1(\alu_shr[14] ),
    .A2(_04693_),
    .B1(_20443_),
    .B2(_04709_),
    .C1(_04712_),
    .X(_02148_));
 sky130_fd_sc_hd__o211a_1 _27072_ (.A1(_04660_),
    .A2(_20446_),
    .B1(_20447_),
    .C1(_04662_),
    .X(_04713_));
 sky130_fd_sc_hd__nor2_1 _27073_ (.A(_04637_),
    .B(_20448_),
    .Y(_04714_));
 sky130_fd_sc_hd__a21o_1 _27074_ (.A1(\alu_shr[15] ),
    .A2(_04633_),
    .B1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__a211o_1 _27075_ (.A1(\alu_shl[15] ),
    .A2(_04658_),
    .B1(_04713_),
    .C1(_04715_),
    .X(_02149_));
 sky130_fd_sc_hd__inv_2 _27076_ (.A(net345),
    .Y(_02363_));
 sky130_fd_sc_hd__a21oi_1 _27077_ (.A1(_02363_),
    .A2(_20776_),
    .B1(_04642_),
    .Y(_04716_));
 sky130_fd_sc_hd__nor2_1 _27078_ (.A(_04637_),
    .B(_20408_),
    .Y(_04717_));
 sky130_fd_sc_hd__a32o_1 _27079_ (.A1(_04668_),
    .A2(net345),
    .A3(_20050_),
    .B1(\alu_shl[16] ),
    .B2(_04652_),
    .X(_04718_));
 sky130_fd_sc_hd__a2111o_1 _27080_ (.A1(_04646_),
    .A2(\alu_shr[16] ),
    .B1(_04716_),
    .C1(_04717_),
    .D1(_04718_),
    .X(_02150_));
 sky130_vsdinv _27081_ (.A(_20395_),
    .Y(_04719_));
 sky130_fd_sc_hd__a22o_1 _27082_ (.A1(\alu_shl[17] ),
    .A2(_04651_),
    .B1(_04670_),
    .B2(\alu_shr[17] ),
    .X(_04720_));
 sky130_fd_sc_hd__a221o_1 _27083_ (.A1(_04719_),
    .A2(_04660_),
    .B1(_20398_),
    .B2(_04648_),
    .C1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__a21o_1 _27084_ (.A1(_20397_),
    .A2(_04669_),
    .B1(_04721_),
    .X(_02151_));
 sky130_fd_sc_hd__or2_1 _27085_ (.A(_20405_),
    .B(_04705_),
    .X(_04722_));
 sky130_vsdinv _27086_ (.A(_20403_),
    .Y(_04723_));
 sky130_fd_sc_hd__a32o_1 _27087_ (.A1(_04694_),
    .A2(_04722_),
    .A3(_04723_),
    .B1(\alu_shl[18] ),
    .B2(_04697_),
    .X(_04724_));
 sky130_fd_sc_hd__a221o_1 _27088_ (.A1(\alu_shr[18] ),
    .A2(_04693_),
    .B1(_20406_),
    .B2(_04709_),
    .C1(_04724_),
    .X(_02152_));
 sky130_fd_sc_hd__or2_1 _27089_ (.A(_20401_),
    .B(_04705_),
    .X(_04725_));
 sky130_vsdinv _27090_ (.A(_20399_),
    .Y(_04726_));
 sky130_fd_sc_hd__a32o_1 _27091_ (.A1(_04694_),
    .A2(_04725_),
    .A3(_04726_),
    .B1(\alu_shl[19] ),
    .B2(_04697_),
    .X(_04727_));
 sky130_fd_sc_hd__a221o_1 _27092_ (.A1(\alu_shr[19] ),
    .A2(_04693_),
    .B1(_20402_),
    .B2(_04709_),
    .C1(_04727_),
    .X(_02153_));
 sky130_fd_sc_hd__o211a_1 _27093_ (.A1(_04659_),
    .A2(_20424_),
    .B1(_20425_),
    .C1(_04662_),
    .X(_04728_));
 sky130_fd_sc_hd__nor2_1 _27094_ (.A(_04637_),
    .B(_20426_),
    .Y(_04729_));
 sky130_fd_sc_hd__a21o_1 _27095_ (.A1(\alu_shl[20] ),
    .A2(_04658_),
    .B1(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__a211o_1 _27096_ (.A1(\alu_shr[20] ),
    .A2(_04646_),
    .B1(_04728_),
    .C1(_04730_),
    .X(_02154_));
 sky130_fd_sc_hd__or2_1 _27097_ (.A(_20416_),
    .B(_04705_),
    .X(_04731_));
 sky130_vsdinv _27098_ (.A(_20414_),
    .Y(_04732_));
 sky130_fd_sc_hd__a32o_1 _27099_ (.A1(_04694_),
    .A2(_04731_),
    .A3(_04732_),
    .B1(\alu_shl[21] ),
    .B2(_04697_),
    .X(_04733_));
 sky130_fd_sc_hd__a221o_1 _27100_ (.A1(\alu_shr[21] ),
    .A2(_04693_),
    .B1(_20417_),
    .B2(_04709_),
    .C1(_04733_),
    .X(_02155_));
 sky130_fd_sc_hd__clkbuf_2 _27101_ (.A(_04645_),
    .X(_04734_));
 sky130_fd_sc_hd__clkbuf_2 _27102_ (.A(_04661_),
    .X(_04735_));
 sky130_fd_sc_hd__or2_1 _27103_ (.A(_20412_),
    .B(_04705_),
    .X(_04736_));
 sky130_vsdinv _27104_ (.A(_20410_),
    .Y(_04737_));
 sky130_fd_sc_hd__clkbuf_2 _27105_ (.A(_04651_),
    .X(_04738_));
 sky130_fd_sc_hd__a32o_1 _27106_ (.A1(_04735_),
    .A2(_04736_),
    .A3(_04737_),
    .B1(\alu_shl[22] ),
    .B2(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__a221o_1 _27107_ (.A1(\alu_shr[22] ),
    .A2(_04734_),
    .B1(_20413_),
    .B2(_04709_),
    .C1(_04739_),
    .X(_02156_));
 sky130_vsdinv _27108_ (.A(_20422_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_1 _27109_ (.A(_20420_),
    .B(_04642_),
    .Y(_04741_));
 sky130_fd_sc_hd__a32o_1 _27110_ (.A1(_04735_),
    .A2(_20421_),
    .A3(_04741_),
    .B1(\alu_shl[23] ),
    .B2(_04738_),
    .X(_04742_));
 sky130_fd_sc_hd__a221o_1 _27111_ (.A1(\alu_shr[23] ),
    .A2(_04734_),
    .B1(_04740_),
    .B2(_04709_),
    .C1(_04742_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_2 _27112_ (.A(_04647_),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_2 _27113_ (.A(_04643_),
    .X(_04744_));
 sky130_fd_sc_hd__or2_1 _27114_ (.A(_20514_),
    .B(_04744_),
    .X(_04745_));
 sky130_vsdinv _27115_ (.A(_20512_),
    .Y(_04746_));
 sky130_fd_sc_hd__a32o_1 _27116_ (.A1(_04735_),
    .A2(_04745_),
    .A3(_04746_),
    .B1(\alu_shl[24] ),
    .B2(_04738_),
    .X(_04747_));
 sky130_fd_sc_hd__a221o_1 _27117_ (.A1(\alu_shr[24] ),
    .A2(_04734_),
    .B1(_20515_),
    .B2(_04743_),
    .C1(_04747_),
    .X(_02158_));
 sky130_fd_sc_hd__or2_1 _27118_ (.A(_20502_),
    .B(_04744_),
    .X(_04748_));
 sky130_vsdinv _27119_ (.A(_20500_),
    .Y(_04749_));
 sky130_fd_sc_hd__a32o_1 _27120_ (.A1(_04735_),
    .A2(_04748_),
    .A3(_04749_),
    .B1(\alu_shl[25] ),
    .B2(_04738_),
    .X(_04750_));
 sky130_fd_sc_hd__a221o_1 _27121_ (.A1(\alu_shr[25] ),
    .A2(_04734_),
    .B1(_20503_),
    .B2(_04743_),
    .C1(_04750_),
    .X(_02159_));
 sky130_fd_sc_hd__or2_1 _27122_ (.A(_20510_),
    .B(_04744_),
    .X(_04751_));
 sky130_vsdinv _27123_ (.A(_20508_),
    .Y(_04752_));
 sky130_fd_sc_hd__a32o_1 _27124_ (.A1(_04735_),
    .A2(_04751_),
    .A3(_04752_),
    .B1(\alu_shl[26] ),
    .B2(_04738_),
    .X(_04753_));
 sky130_fd_sc_hd__a221o_1 _27125_ (.A1(\alu_shr[26] ),
    .A2(_04734_),
    .B1(_20511_),
    .B2(_04743_),
    .C1(_04753_),
    .X(_02160_));
 sky130_fd_sc_hd__or2_1 _27126_ (.A(_20523_),
    .B(_04744_),
    .X(_04754_));
 sky130_vsdinv _27127_ (.A(_20521_),
    .Y(_04755_));
 sky130_fd_sc_hd__a32o_1 _27128_ (.A1(_04735_),
    .A2(_04754_),
    .A3(_04755_),
    .B1(\alu_shl[27] ),
    .B2(_04738_),
    .X(_04756_));
 sky130_fd_sc_hd__a221o_1 _27129_ (.A1(\alu_shr[27] ),
    .A2(_04734_),
    .B1(_20524_),
    .B2(_04743_),
    .C1(_04756_),
    .X(_02161_));
 sky130_fd_sc_hd__or2_1 _27130_ (.A(_20506_),
    .B(_04744_),
    .X(_04757_));
 sky130_vsdinv _27131_ (.A(_20504_),
    .Y(_04758_));
 sky130_fd_sc_hd__a32o_1 _27132_ (.A1(_04661_),
    .A2(_04757_),
    .A3(_04758_),
    .B1(\alu_shl[28] ),
    .B2(_04657_),
    .X(_04759_));
 sky130_fd_sc_hd__a221o_1 _27133_ (.A1(\alu_shr[28] ),
    .A2(_04633_),
    .B1(_20507_),
    .B2(_04743_),
    .C1(_04759_),
    .X(_02162_));
 sky130_vsdinv _27134_ (.A(_20517_),
    .Y(_04760_));
 sky130_fd_sc_hd__a22o_1 _27135_ (.A1(_04658_),
    .A2(\alu_shl[29] ),
    .B1(_20519_),
    .B2(_04668_),
    .X(_04761_));
 sky130_fd_sc_hd__a22o_1 _27136_ (.A1(_20520_),
    .A2(_04648_),
    .B1(_04633_),
    .B2(\alu_shr[29] ),
    .X(_04762_));
 sky130_fd_sc_hd__a211o_1 _27137_ (.A1(_04760_),
    .A2(_04667_),
    .B1(_04761_),
    .C1(_04762_),
    .X(_02163_));
 sky130_vsdinv _27138_ (.A(_20528_),
    .Y(_04763_));
 sky130_fd_sc_hd__a22o_1 _27139_ (.A1(\alu_shl[30] ),
    .A2(_04651_),
    .B1(_04670_),
    .B2(\alu_shr[30] ),
    .X(_04764_));
 sky130_fd_sc_hd__a221o_1 _27140_ (.A1(_04763_),
    .A2(_04660_),
    .B1(_20531_),
    .B2(_04648_),
    .C1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a21o_1 _27141_ (.A1(_20530_),
    .A2(_04669_),
    .B1(_04765_),
    .X(_02164_));
 sky130_fd_sc_hd__or2_1 _27142_ (.A(_20526_),
    .B(_04744_),
    .X(_04766_));
 sky130_vsdinv _27143_ (.A(_20525_),
    .Y(_04767_));
 sky130_fd_sc_hd__a32o_1 _27144_ (.A1(_04661_),
    .A2(_04766_),
    .A3(_04767_),
    .B1(\alu_shl[31] ),
    .B2(_04657_),
    .X(_04768_));
 sky130_fd_sc_hd__a221o_1 _27145_ (.A1(\alu_shr[31] ),
    .A2(_04633_),
    .B1(_20527_),
    .B2(_04743_),
    .C1(_04768_),
    .X(_02165_));
 sky130_fd_sc_hd__and3_1 _27146_ (.A(_00289_),
    .B(_18525_),
    .C(_20551_),
    .X(_02166_));
 sky130_fd_sc_hd__buf_2 _27147_ (.A(\mem_wordsize[1] ),
    .X(_04769_));
 sky130_fd_sc_hd__a22o_1 _27148_ (.A1(net368),
    .A2(_04166_),
    .B1(_19677_),
    .B2(_04769_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_1 _27149_ (.A1(_19668_),
    .A2(_04166_),
    .B1(_19676_),
    .B2(_04769_),
    .X(_02168_));
 sky130_fd_sc_hd__buf_2 _27150_ (.A(_04094_),
    .X(_04770_));
 sky130_fd_sc_hd__a22o_1 _27151_ (.A1(net339),
    .A2(_04770_),
    .B1(_19675_),
    .B2(_04769_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _27152_ (.A1(_19667_),
    .A2(_04770_),
    .B1(_20311_),
    .B2(_04769_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _27153_ (.A1(net341),
    .A2(_04770_),
    .B1(_19673_),
    .B2(_04769_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_1 _27154_ (.A1(_19666_),
    .A2(_04770_),
    .B1(_19672_),
    .B2(_04769_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_1 _27155_ (.A1(net343),
    .A2(_04770_),
    .B1(_19671_),
    .B2(\mem_wordsize[1] ),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_1 _27156_ (.A1(_19664_),
    .A2(_04770_),
    .B1(_19670_),
    .B2(\mem_wordsize[1] ),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_1 _27157_ (.A(_20392_),
    .B(_04466_),
    .Y(_02175_));
 sky130_fd_sc_hd__clkbuf_2 _27158_ (.A(_04093_),
    .X(_04771_));
 sky130_fd_sc_hd__nor2_1 _27159_ (.A(_02318_),
    .B(_04771_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _27160_ (.A(_02321_),
    .B(_04771_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _27161_ (.A(_02324_),
    .B(_04771_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _27162_ (.A(_02327_),
    .B(_04771_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _27163_ (.A(_02330_),
    .B(_04771_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _27164_ (.A(_02333_),
    .B(_04771_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _27165_ (.A(_02336_),
    .B(_04093_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_8 _27166_ (.A(_20555_),
    .B(net511),
    .Y(_02183_));
 sky130_fd_sc_hd__or2_1 _27167_ (.A(\irq_pending[3] ),
    .B(net26),
    .X(_02214_));
 sky130_fd_sc_hd__and2_1 _27168_ (.A(_02214_),
    .B(\irq_mask[3] ),
    .X(_02215_));
 sky130_vsdinv _27169_ (.A(_01700_),
    .Y(_02217_));
 sky130_fd_sc_hd__or2_1 _27170_ (.A(\irq_pending[4] ),
    .B(net27),
    .X(_02218_));
 sky130_fd_sc_hd__and2_1 _27171_ (.A(_02218_),
    .B(\irq_mask[4] ),
    .X(_02219_));
 sky130_fd_sc_hd__or2_1 _27172_ (.A(\irq_pending[5] ),
    .B(net28),
    .X(_02221_));
 sky130_fd_sc_hd__and2_1 _27173_ (.A(_02221_),
    .B(\irq_mask[5] ),
    .X(_02222_));
 sky130_fd_sc_hd__or2_1 _27174_ (.A(\irq_pending[6] ),
    .B(net29),
    .X(_02224_));
 sky130_fd_sc_hd__and2_1 _27175_ (.A(_02224_),
    .B(\irq_mask[6] ),
    .X(_02225_));
 sky130_fd_sc_hd__or2_1 _27176_ (.A(\irq_pending[7] ),
    .B(net529),
    .X(_02227_));
 sky130_fd_sc_hd__and2_1 _27177_ (.A(_02227_),
    .B(\irq_mask[7] ),
    .X(_02228_));
 sky130_fd_sc_hd__or2_1 _27178_ (.A(\irq_pending[8] ),
    .B(net31),
    .X(_02230_));
 sky130_fd_sc_hd__and2_1 _27179_ (.A(_02230_),
    .B(\irq_mask[8] ),
    .X(_02231_));
 sky130_fd_sc_hd__or2_1 _27180_ (.A(\irq_pending[9] ),
    .B(net32),
    .X(_02233_));
 sky130_fd_sc_hd__and2_1 _27181_ (.A(_02233_),
    .B(\irq_mask[9] ),
    .X(_02234_));
 sky130_fd_sc_hd__or2_1 _27182_ (.A(\irq_pending[10] ),
    .B(net532),
    .X(_02236_));
 sky130_fd_sc_hd__and2_1 _27183_ (.A(_02236_),
    .B(\irq_mask[10] ),
    .X(_02237_));
 sky130_fd_sc_hd__or2_1 _27184_ (.A(\irq_pending[11] ),
    .B(net3),
    .X(_02239_));
 sky130_fd_sc_hd__and2_1 _27185_ (.A(_02239_),
    .B(\irq_mask[11] ),
    .X(_02240_));
 sky130_fd_sc_hd__or2_1 _27186_ (.A(\irq_pending[12] ),
    .B(net4),
    .X(_02242_));
 sky130_fd_sc_hd__and2_1 _27187_ (.A(_02242_),
    .B(\irq_mask[12] ),
    .X(_02243_));
 sky130_fd_sc_hd__or2_1 _27188_ (.A(\irq_pending[13] ),
    .B(net5),
    .X(_02245_));
 sky130_fd_sc_hd__and2_1 _27189_ (.A(_02245_),
    .B(\irq_mask[13] ),
    .X(_02246_));
 sky130_fd_sc_hd__or2_1 _27190_ (.A(\irq_pending[14] ),
    .B(net6),
    .X(_02248_));
 sky130_fd_sc_hd__and2_1 _27191_ (.A(_02248_),
    .B(\irq_mask[14] ),
    .X(_02249_));
 sky130_fd_sc_hd__or2_1 _27192_ (.A(\irq_pending[15] ),
    .B(net520),
    .X(_02251_));
 sky130_fd_sc_hd__and2_1 _27193_ (.A(_02251_),
    .B(\irq_mask[15] ),
    .X(_02252_));
 sky130_fd_sc_hd__or2_1 _27194_ (.A(\irq_pending[16] ),
    .B(net8),
    .X(_02254_));
 sky130_fd_sc_hd__and2_1 _27195_ (.A(_02254_),
    .B(\irq_mask[16] ),
    .X(_02255_));
 sky130_fd_sc_hd__or2_1 _27196_ (.A(\irq_pending[17] ),
    .B(net9),
    .X(_02257_));
 sky130_fd_sc_hd__and2_1 _27197_ (.A(_02257_),
    .B(\irq_mask[17] ),
    .X(_02258_));
 sky130_fd_sc_hd__or2_1 _27198_ (.A(\irq_pending[18] ),
    .B(net10),
    .X(_02260_));
 sky130_fd_sc_hd__and2_1 _27199_ (.A(_02260_),
    .B(\irq_mask[18] ),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _27200_ (.A(\irq_pending[19] ),
    .B(net11),
    .X(_02263_));
 sky130_fd_sc_hd__and2_1 _27201_ (.A(_02263_),
    .B(\irq_mask[19] ),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _27202_ (.A(\irq_pending[20] ),
    .B(net533),
    .X(_02266_));
 sky130_fd_sc_hd__and2_1 _27203_ (.A(_02266_),
    .B(\irq_mask[20] ),
    .X(_02267_));
 sky130_fd_sc_hd__or2_1 _27204_ (.A(\irq_pending[21] ),
    .B(net14),
    .X(_02269_));
 sky130_fd_sc_hd__and2_1 _27205_ (.A(_02269_),
    .B(\irq_mask[21] ),
    .X(_02270_));
 sky130_fd_sc_hd__or2_1 _27206_ (.A(\irq_pending[22] ),
    .B(net15),
    .X(_02272_));
 sky130_fd_sc_hd__and2_1 _27207_ (.A(_02272_),
    .B(\irq_mask[22] ),
    .X(_02273_));
 sky130_fd_sc_hd__or2_1 _27208_ (.A(\irq_pending[23] ),
    .B(net16),
    .X(_02275_));
 sky130_fd_sc_hd__and2_1 _27209_ (.A(_02275_),
    .B(\irq_mask[23] ),
    .X(_02276_));
 sky130_fd_sc_hd__or2_1 _27210_ (.A(\irq_pending[24] ),
    .B(net17),
    .X(_02278_));
 sky130_fd_sc_hd__and2_1 _27211_ (.A(_02278_),
    .B(\irq_mask[24] ),
    .X(_02279_));
 sky130_fd_sc_hd__or2_1 _27212_ (.A(\irq_pending[25] ),
    .B(net18),
    .X(_02281_));
 sky130_fd_sc_hd__and2_1 _27213_ (.A(_02281_),
    .B(\irq_mask[25] ),
    .X(_02282_));
 sky130_fd_sc_hd__or2_1 _27214_ (.A(\irq_pending[26] ),
    .B(net19),
    .X(_02284_));
 sky130_fd_sc_hd__and2_1 _27215_ (.A(_02284_),
    .B(\irq_mask[26] ),
    .X(_02285_));
 sky130_fd_sc_hd__or2_1 _27216_ (.A(\irq_pending[27] ),
    .B(net531),
    .X(_02287_));
 sky130_fd_sc_hd__and2_1 _27217_ (.A(_02287_),
    .B(\irq_mask[27] ),
    .X(_02288_));
 sky130_fd_sc_hd__or2_1 _27218_ (.A(\irq_pending[28] ),
    .B(net530),
    .X(_02290_));
 sky130_fd_sc_hd__and2_1 _27219_ (.A(_02290_),
    .B(\irq_mask[28] ),
    .X(_02291_));
 sky130_fd_sc_hd__or2_1 _27220_ (.A(\irq_pending[29] ),
    .B(net22),
    .X(_02293_));
 sky130_fd_sc_hd__and2_1 _27221_ (.A(_02293_),
    .B(\irq_mask[29] ),
    .X(_02294_));
 sky130_fd_sc_hd__or2_1 _27222_ (.A(\irq_pending[30] ),
    .B(net24),
    .X(_02296_));
 sky130_fd_sc_hd__and2_1 _27223_ (.A(_02296_),
    .B(\irq_mask[30] ),
    .X(_02297_));
 sky130_fd_sc_hd__or2_1 _27224_ (.A(\irq_pending[31] ),
    .B(net25),
    .X(_02299_));
 sky130_fd_sc_hd__and2_1 _27225_ (.A(_02299_),
    .B(\irq_mask[31] ),
    .X(_02300_));
 sky130_fd_sc_hd__nor2_1 _27226_ (.A(\timer[27] ),
    .B(\timer[26] ),
    .Y(_04772_));
 sky130_fd_sc_hd__and3b_1 _27227_ (.A_N(_20556_),
    .B(_20587_),
    .C(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__or2_1 _27228_ (.A(\timer[11] ),
    .B(\timer[10] ),
    .X(_04774_));
 sky130_fd_sc_hd__or2_1 _27229_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .X(_04775_));
 sky130_fd_sc_hd__or4_4 _27230_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(\timer[7] ),
    .D(\timer[6] ),
    .X(_04776_));
 sky130_fd_sc_hd__nor3_2 _27231_ (.A(_04774_),
    .B(_04775_),
    .C(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__and4_1 _27232_ (.A(_20580_),
    .B(_04515_),
    .C(_04504_),
    .D(_20583_),
    .X(_04778_));
 sky130_fd_sc_hd__and4_1 _27233_ (.A(_04127_),
    .B(_04317_),
    .C(_20574_),
    .D(\timer[0] ),
    .X(_04779_));
 sky130_fd_sc_hd__and3_1 _27234_ (.A(_04779_),
    .B(_20557_),
    .C(_20568_),
    .X(_04780_));
 sky130_fd_sc_hd__a41o_1 _27235_ (.A1(_04773_),
    .A2(_04777_),
    .A3(_04778_),
    .A4(_04780_),
    .B1(\irq_pending[0] ),
    .X(_02302_));
 sky130_fd_sc_hd__or2_1 _27236_ (.A(_02303_),
    .B(net1),
    .X(_02304_));
 sky130_fd_sc_hd__and2_1 _27237_ (.A(_02304_),
    .B(\irq_mask[0] ),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_1 _27238_ (.A(\irq_pending[2] ),
    .B(net23),
    .Y(_02307_));
 sky130_fd_sc_hd__or2_1 _27239_ (.A(_18595_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__nor2_1 _27240_ (.A(_02310_),
    .B(_19506_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_1 _27241_ (.A(_20338_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__or2_1 _27242_ (.A(_02313_),
    .B(_20338_),
    .X(_02314_));
 sky130_fd_sc_hd__or2_1 _27243_ (.A(_02316_),
    .B(_20338_),
    .X(_02317_));
 sky130_fd_sc_hd__or3_1 _27244_ (.A(_02387_),
    .B(net322),
    .C(_20503_),
    .X(_04781_));
 sky130_fd_sc_hd__nand2_1 _27245_ (.A(_20501_),
    .B(_19659_),
    .Y(_04782_));
 sky130_fd_sc_hd__a21o_1 _27246_ (.A1(_04781_),
    .A2(_04782_),
    .B1(_20511_),
    .X(_04783_));
 sky130_fd_sc_hd__nand2_1 _27247_ (.A(_20509_),
    .B(_19657_),
    .Y(_04784_));
 sky130_fd_sc_hd__a21o_1 _27248_ (.A1(_04783_),
    .A2(_04784_),
    .B1(_20524_),
    .X(_04785_));
 sky130_fd_sc_hd__nand2_1 _27249_ (.A(_20522_),
    .B(_19656_),
    .Y(_04786_));
 sky130_fd_sc_hd__a211o_1 _27250_ (.A1(_04785_),
    .A2(_04786_),
    .B1(_20507_),
    .C1(_20520_),
    .X(_04787_));
 sky130_fd_sc_hd__nand2_1 _27251_ (.A(_20518_),
    .B(_19655_),
    .Y(_04788_));
 sky130_fd_sc_hd__or3_1 _27252_ (.A(_02399_),
    .B(_20038_),
    .C(_20520_),
    .X(_04789_));
 sky130_fd_sc_hd__a311o_1 _27253_ (.A1(_04787_),
    .A2(_04788_),
    .A3(_04789_),
    .B1(_20527_),
    .C1(_20531_),
    .X(_04790_));
 sky130_vsdinv _27254_ (.A(_20321_),
    .Y(_04791_));
 sky130_fd_sc_hd__nor2_2 _27255_ (.A(_20322_),
    .B(_04791_),
    .Y(_00049_));
 sky130_fd_sc_hd__o21a_1 _27256_ (.A1(_20320_),
    .A2(_00048_),
    .B1(_20063_),
    .X(_04792_));
 sky130_fd_sc_hd__or3b_2 _27257_ (.A(_00049_),
    .B(_04792_),
    .C_N(_20485_),
    .X(_04793_));
 sky130_fd_sc_hd__nand2_1 _27258_ (.A(_20478_),
    .B(_19674_),
    .Y(_04794_));
 sky130_fd_sc_hd__or3_1 _27259_ (.A(_20319_),
    .B(_20062_),
    .C(_20480_),
    .X(_04795_));
 sky130_fd_sc_hd__a311o_1 _27260_ (.A1(_04793_),
    .A2(_04794_),
    .A3(_04795_),
    .B1(_20471_),
    .C1(_20490_),
    .X(_04796_));
 sky130_fd_sc_hd__nand2_1 _27261_ (.A(_20469_),
    .B(_19672_),
    .Y(_04797_));
 sky130_fd_sc_hd__or3_1 _27262_ (.A(_20310_),
    .B(_20060_),
    .C(_20471_),
    .X(_04798_));
 sky130_fd_sc_hd__a31o_1 _27263_ (.A1(_04796_),
    .A2(_04797_),
    .A3(_04798_),
    .B1(_20476_),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_1 _27264_ (.A(_20472_),
    .B(_19671_),
    .Y(_04800_));
 sky130_fd_sc_hd__a21bo_1 _27265_ (.A1(_04799_),
    .A2(_04800_),
    .B1_N(_20497_),
    .X(_04801_));
 sky130_fd_sc_hd__nand2_1 _27266_ (.A(_20703_),
    .B(net229),
    .Y(_04802_));
 sky130_fd_sc_hd__a21o_1 _27267_ (.A1(_04801_),
    .A2(_04802_),
    .B1(_20467_),
    .X(_04803_));
 sky130_fd_sc_hd__nand2_1 _27268_ (.A(_20452_),
    .B(_19667_),
    .Y(_04804_));
 sky130_fd_sc_hd__or3_2 _27269_ (.A(_02339_),
    .B(_20056_),
    .C(_20458_),
    .X(_04805_));
 sky130_fd_sc_hd__nand2_1 _27270_ (.A(_20456_),
    .B(_19668_),
    .Y(_04806_));
 sky130_fd_sc_hd__a21o_1 _27271_ (.A1(_04805_),
    .A2(_04806_),
    .B1(_20466_),
    .X(_04807_));
 sky130_fd_sc_hd__nand2_1 _27272_ (.A(_20464_),
    .B(net339),
    .Y(_04808_));
 sky130_fd_sc_hd__a21o_1 _27273_ (.A1(_04807_),
    .A2(_04808_),
    .B1(_20454_),
    .X(_04809_));
 sky130_fd_sc_hd__a31o_1 _27274_ (.A1(_04803_),
    .A2(_04804_),
    .A3(_04809_),
    .B1(_20450_),
    .X(_04810_));
 sky130_fd_sc_hd__nand2_1 _27275_ (.A(_20445_),
    .B(_19664_),
    .Y(_04811_));
 sky130_fd_sc_hd__nor2_1 _27276_ (.A(_20051_),
    .B(_02357_),
    .Y(_04812_));
 sky130_fd_sc_hd__or3_1 _27277_ (.A(_02351_),
    .B(_20053_),
    .C(_20433_),
    .X(_04813_));
 sky130_fd_sc_hd__nand2_1 _27278_ (.A(_20431_),
    .B(_19666_),
    .Y(_04814_));
 sky130_fd_sc_hd__a21oi_1 _27279_ (.A1(_04813_),
    .A2(_04814_),
    .B1(_20443_),
    .Y(_04815_));
 sky130_fd_sc_hd__o21ai_1 _27280_ (.A1(_04812_),
    .A2(_04815_),
    .B1(_20448_),
    .Y(_04816_));
 sky130_fd_sc_hd__a31o_1 _27281_ (.A1(_04810_),
    .A2(_04811_),
    .A3(_04816_),
    .B1(_20429_),
    .X(_04817_));
 sky130_fd_sc_hd__nor2_1 _27282_ (.A(_20044_),
    .B(_02381_),
    .Y(_04818_));
 sky130_fd_sc_hd__or3_1 _27283_ (.A(_02375_),
    .B(_20046_),
    .C(_20417_),
    .X(_04819_));
 sky130_fd_sc_hd__nand2_1 _27284_ (.A(_20415_),
    .B(_19660_),
    .Y(_04820_));
 sky130_fd_sc_hd__a21oi_1 _27285_ (.A1(_04819_),
    .A2(_04820_),
    .B1(_20413_),
    .Y(_04821_));
 sky130_fd_sc_hd__o21ai_1 _27286_ (.A1(_04818_),
    .A2(_04821_),
    .B1(_20422_),
    .Y(_04822_));
 sky130_fd_sc_hd__or3_1 _27287_ (.A(_02363_),
    .B(_20050_),
    .C(_20398_),
    .X(_04823_));
 sky130_fd_sc_hd__nand2_1 _27288_ (.A(_20396_),
    .B(_19663_),
    .Y(_04824_));
 sky130_fd_sc_hd__a21o_1 _27289_ (.A1(_04823_),
    .A2(_04824_),
    .B1(_20406_),
    .X(_04825_));
 sky130_fd_sc_hd__nand2_1 _27290_ (.A(_20404_),
    .B(_19662_),
    .Y(_04826_));
 sky130_fd_sc_hd__a21o_1 _27291_ (.A1(_04825_),
    .A2(_04826_),
    .B1(_20402_),
    .X(_04827_));
 sky130_fd_sc_hd__nand2_1 _27292_ (.A(_20400_),
    .B(net348),
    .Y(_04828_));
 sky130_fd_sc_hd__a21o_1 _27293_ (.A1(_04827_),
    .A2(_04828_),
    .B1(_20428_),
    .X(_04829_));
 sky130_fd_sc_hd__o211a_1 _27294_ (.A1(_02384_),
    .A2(_20043_),
    .B1(_04822_),
    .C1(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__a21bo_1 _27295_ (.A1(_04817_),
    .A2(_04830_),
    .B1_N(_20533_),
    .X(_04831_));
 sky130_fd_sc_hd__o311a_4 _27296_ (.A1(_02405_),
    .A2(_20036_),
    .A3(_20527_),
    .B1(_04790_),
    .C1(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__nor2_2 _27297_ (.A(net330),
    .B(_18690_),
    .Y(_04833_));
 sky130_vsdinv _27298_ (.A(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__a21oi_1 _27299_ (.A1(_04832_),
    .A2(_04834_),
    .B1(_00000_),
    .Y(_00002_));
 sky130_vsdinv _27300_ (.A(_20527_),
    .Y(_04835_));
 sky130_fd_sc_hd__a211oi_4 _27301_ (.A1(_04832_),
    .A2(_04835_),
    .B1(_00000_),
    .C1(_04833_),
    .Y(_00001_));
 sky130_vsdinv _27302_ (.A(\pcpi_mul.rs2[0] ),
    .Y(_04836_));
 sky130_fd_sc_hd__clkbuf_2 _27303_ (.A(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__buf_6 _27304_ (.A(\pcpi_mul.rs1[0] ),
    .X(_04838_));
 sky130_fd_sc_hd__clkinv_8 _27305_ (.A(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__clkbuf_2 _27306_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__buf_8 _27307_ (.A(net449),
    .X(_04841_));
 sky130_fd_sc_hd__nor2_2 _27308_ (.A(net470),
    .B(_04841_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _27309_ (.A(_19676_),
    .B(_19677_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand2_1 _27310_ (.A(_04791_),
    .B(_04842_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _27311_ (.A(net317),
    .B(_02320_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_1 _27312_ (.A(net317),
    .B(_02320_),
    .Y(_04844_));
 sky130_fd_sc_hd__or2b_1 _27313_ (.A(_04843_),
    .B_N(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__xor2_1 _27314_ (.A(_20393_),
    .B(_04845_),
    .X(_02602_));
 sky130_fd_sc_hd__nor2_1 _27315_ (.A(_19675_),
    .B(_04791_),
    .Y(_04846_));
 sky130_vsdinv _27316_ (.A(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _27317_ (.A(_04791_),
    .B(_19675_),
    .Y(_04848_));
 sky130_fd_sc_hd__nand2_1 _27318_ (.A(_04847_),
    .B(_04848_),
    .Y(_02322_));
 sky130_fd_sc_hd__o21ai_2 _27319_ (.A1(_04843_),
    .A2(_20393_),
    .B1(_04844_),
    .Y(_04849_));
 sky130_vsdinv _27320_ (.A(_02323_),
    .Y(_04850_));
 sky130_fd_sc_hd__nor2_2 _27321_ (.A(_20482_),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand2_2 _27322_ (.A(_20482_),
    .B(_04850_),
    .Y(_04852_));
 sky130_fd_sc_hd__and2b_1 _27323_ (.A_N(_04851_),
    .B(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__xor2_1 _27324_ (.A(_04849_),
    .B(_04853_),
    .X(_02613_));
 sky130_fd_sc_hd__nand2_1 _27325_ (.A(_04847_),
    .B(_20311_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _27326_ (.A(_04854_),
    .B(_20324_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_1 _27327_ (.A(_20061_),
    .B(_02326_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _27328_ (.A(_20061_),
    .B(_02326_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2b_1 _27329_ (.A(_04855_),
    .B_N(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__a21oi_4 _27330_ (.A1(_04849_),
    .A2(_04852_),
    .B1(_04851_),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_1 _27331_ (.A(_04857_),
    .B(_04858_),
    .X(_02616_));
 sky130_fd_sc_hd__nand2_1 _27332_ (.A(_20324_),
    .B(_19673_),
    .Y(_04859_));
 sky130_fd_sc_hd__nand2_1 _27333_ (.A(_20326_),
    .B(_04859_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_1 _27334_ (.A(_20060_),
    .B(_02329_),
    .Y(_04860_));
 sky130_fd_sc_hd__and2_1 _27335_ (.A(_20060_),
    .B(_02329_),
    .X(_04861_));
 sky130_fd_sc_hd__nor2_1 _27336_ (.A(_04860_),
    .B(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__o21ai_2 _27337_ (.A1(_04855_),
    .A2(_04858_),
    .B1(_04856_),
    .Y(_04863_));
 sky130_fd_sc_hd__xor2_1 _27338_ (.A(_04862_),
    .B(_04863_),
    .X(_02617_));
 sky130_fd_sc_hd__nand2_1 _27339_ (.A(_20326_),
    .B(_19672_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_1 _27340_ (.A(_20325_),
    .B(_02330_),
    .Y(_04865_));
 sky130_fd_sc_hd__nand2_1 _27341_ (.A(_04864_),
    .B(_04865_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _27342_ (.A(_20059_),
    .B(_02332_),
    .Y(_04866_));
 sky130_fd_sc_hd__nand2_1 _27343_ (.A(_20059_),
    .B(_02332_),
    .Y(_04867_));
 sky130_fd_sc_hd__or2b_1 _27344_ (.A(_04866_),
    .B_N(_04867_),
    .X(_04868_));
 sky130_vsdinv _27345_ (.A(_04860_),
    .Y(_04869_));
 sky130_fd_sc_hd__a21oi_4 _27346_ (.A1(_04863_),
    .A2(_04869_),
    .B1(_04861_),
    .Y(_04870_));
 sky130_fd_sc_hd__xor2_1 _27347_ (.A(_04868_),
    .B(_04870_),
    .X(_02618_));
 sky130_fd_sc_hd__or2_1 _27348_ (.A(net228),
    .B(_04865_),
    .X(_04871_));
 sky130_fd_sc_hd__nand2_1 _27349_ (.A(_04865_),
    .B(_19671_),
    .Y(_04872_));
 sky130_fd_sc_hd__nand2_1 _27350_ (.A(_04871_),
    .B(_04872_),
    .Y(_02334_));
 sky130_fd_sc_hd__or2_1 _27351_ (.A(net334),
    .B(_02335_),
    .X(_04873_));
 sky130_fd_sc_hd__nand2_1 _27352_ (.A(net334),
    .B(_02335_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_1 _27353_ (.A(_04873_),
    .B(_04874_),
    .Y(_04875_));
 sky130_vsdinv _27354_ (.A(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__o21ai_2 _27355_ (.A1(_04866_),
    .A2(_04870_),
    .B1(_04867_),
    .Y(_04877_));
 sky130_fd_sc_hd__or2_1 _27356_ (.A(_04876_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _27357_ (.A(_04877_),
    .B(_04876_),
    .Y(_04879_));
 sky130_fd_sc_hd__and2_1 _27358_ (.A(_04878_),
    .B(_04879_),
    .X(_02619_));
 sky130_fd_sc_hd__nor2_2 _27359_ (.A(net229),
    .B(_04871_),
    .Y(_04880_));
 sky130_fd_sc_hd__and2_1 _27360_ (.A(_04871_),
    .B(_19670_),
    .X(_04881_));
 sky130_fd_sc_hd__or2_1 _27361_ (.A(_04880_),
    .B(_04881_),
    .X(_02337_));
 sky130_fd_sc_hd__nor2_1 _27362_ (.A(_20057_),
    .B(_02338_),
    .Y(_04882_));
 sky130_vsdinv _27363_ (.A(_02338_),
    .Y(_04883_));
 sky130_fd_sc_hd__nor2_1 _27364_ (.A(_20703_),
    .B(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nor2_1 _27365_ (.A(_04882_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _27366_ (.A(_04879_),
    .B(_04874_),
    .Y(_04886_));
 sky130_fd_sc_hd__xor2_1 _27367_ (.A(_04885_),
    .B(_04886_),
    .X(_02620_));
 sky130_fd_sc_hd__or2_1 _27368_ (.A(_02339_),
    .B(_04880_),
    .X(_04887_));
 sky130_fd_sc_hd__nand2_1 _27369_ (.A(_04880_),
    .B(_02339_),
    .Y(_04888_));
 sky130_fd_sc_hd__nand2_1 _27370_ (.A(_04887_),
    .B(_04888_),
    .Y(_02340_));
 sky130_fd_sc_hd__or2_1 _27371_ (.A(_20056_),
    .B(_02341_),
    .X(_04889_));
 sky130_fd_sc_hd__nand2_1 _27372_ (.A(_20056_),
    .B(_02341_),
    .Y(_04890_));
 sky130_fd_sc_hd__and2_1 _27373_ (.A(_04889_),
    .B(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__and3_1 _27374_ (.A(_04885_),
    .B(_04874_),
    .C(_04873_),
    .X(_04892_));
 sky130_fd_sc_hd__o21ba_1 _27375_ (.A1(_04874_),
    .A2(_04882_),
    .B1_N(_04884_),
    .X(_04893_));
 sky130_fd_sc_hd__a21boi_1 _27376_ (.A1(_04877_),
    .A2(_04892_),
    .B1_N(_04893_),
    .Y(_04894_));
 sky130_vsdinv _27377_ (.A(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__or2_1 _27378_ (.A(_04891_),
    .B(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__nand2_1 _27379_ (.A(_04895_),
    .B(_04891_),
    .Y(_04897_));
 sky130_fd_sc_hd__and2_1 _27380_ (.A(_04896_),
    .B(_04897_),
    .X(_02621_));
 sky130_fd_sc_hd__nor2_1 _27381_ (.A(net369),
    .B(_04888_),
    .Y(_04898_));
 sky130_fd_sc_hd__and2_1 _27382_ (.A(_04888_),
    .B(_19668_),
    .X(_04899_));
 sky130_fd_sc_hd__or2_1 _27383_ (.A(_04898_),
    .B(_04899_),
    .X(_02343_));
 sky130_fd_sc_hd__nor2_1 _27384_ (.A(_20055_),
    .B(_02344_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _27385_ (.A(_20055_),
    .B(_02344_),
    .Y(_04901_));
 sky130_fd_sc_hd__and2b_1 _27386_ (.A_N(_04900_),
    .B(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__nand2_1 _27387_ (.A(_04897_),
    .B(_04890_),
    .Y(_04903_));
 sky130_fd_sc_hd__xor2_1 _27388_ (.A(_04902_),
    .B(_04903_),
    .X(_02622_));
 sky130_fd_sc_hd__or2_1 _27389_ (.A(_02345_),
    .B(_04898_),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _27390_ (.A(_04898_),
    .B(_02345_),
    .Y(_04905_));
 sky130_fd_sc_hd__nand2_1 _27391_ (.A(_04904_),
    .B(_04905_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _27392_ (.A(_20054_),
    .B(_02347_),
    .Y(_04906_));
 sky130_fd_sc_hd__nand2_1 _27393_ (.A(_20054_),
    .B(_02347_),
    .Y(_04907_));
 sky130_vsdinv _27394_ (.A(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__nor2_2 _27395_ (.A(_04906_),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand2_1 _27396_ (.A(_04891_),
    .B(_04902_),
    .Y(_04910_));
 sky130_fd_sc_hd__o21a_1 _27397_ (.A1(_04890_),
    .A2(_04900_),
    .B1(_04901_),
    .X(_04911_));
 sky130_fd_sc_hd__o21ai_1 _27398_ (.A1(_04910_),
    .A2(_04894_),
    .B1(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__or2_1 _27399_ (.A(_04909_),
    .B(_04912_),
    .X(_04913_));
 sky130_vsdinv _27400_ (.A(_04911_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _27401_ (.A(_04877_),
    .B(_04892_),
    .Y(_04915_));
 sky130_fd_sc_hd__a21oi_2 _27402_ (.A1(_04915_),
    .A2(_04893_),
    .B1(_04910_),
    .Y(_04916_));
 sky130_fd_sc_hd__o21ai_2 _27403_ (.A1(_04914_),
    .A2(_04916_),
    .B1(_04909_),
    .Y(_04917_));
 sky130_fd_sc_hd__and2_1 _27404_ (.A(_04913_),
    .B(_04917_),
    .X(_02592_));
 sky130_fd_sc_hd__nor2_1 _27405_ (.A(net340),
    .B(_04905_),
    .Y(_04918_));
 sky130_fd_sc_hd__and2_1 _27406_ (.A(_04905_),
    .B(_19667_),
    .X(_04919_));
 sky130_fd_sc_hd__or2_1 _27407_ (.A(_04918_),
    .B(_04919_),
    .X(_02349_));
 sky130_vsdinv _27408_ (.A(_02350_),
    .Y(_04920_));
 sky130_fd_sc_hd__nor2_2 _27409_ (.A(_20452_),
    .B(_04920_),
    .Y(_04921_));
 sky130_vsdinv _27410_ (.A(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_1 _27411_ (.A(_20452_),
    .B(_04920_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _27412_ (.A(_04922_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__a21oi_2 _27413_ (.A1(_04917_),
    .A2(_04907_),
    .B1(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__and3_1 _27414_ (.A(_04917_),
    .B(_04907_),
    .C(_04924_),
    .X(_04926_));
 sky130_fd_sc_hd__nor2_1 _27415_ (.A(_04925_),
    .B(_04926_),
    .Y(_02593_));
 sky130_fd_sc_hd__or2_1 _27416_ (.A(_02351_),
    .B(_04918_),
    .X(_04927_));
 sky130_fd_sc_hd__nand2_1 _27417_ (.A(_04918_),
    .B(_02351_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _27418_ (.A(_04927_),
    .B(_04928_),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_1 _27419_ (.A(_20053_),
    .B(_02353_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _27420_ (.A(_20053_),
    .B(_02353_),
    .Y(_04930_));
 sky130_vsdinv _27421_ (.A(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__nor2_2 _27422_ (.A(_04929_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__a21oi_1 _27423_ (.A1(_04912_),
    .A2(_04909_),
    .B1(_04908_),
    .Y(_04933_));
 sky130_fd_sc_hd__o21ai_1 _27424_ (.A1(_04924_),
    .A2(_04933_),
    .B1(_04922_),
    .Y(_04934_));
 sky130_fd_sc_hd__or2_1 _27425_ (.A(_04932_),
    .B(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__o21ai_2 _27426_ (.A1(_04921_),
    .A2(_04925_),
    .B1(_04932_),
    .Y(_04936_));
 sky130_fd_sc_hd__and2_1 _27427_ (.A(_04935_),
    .B(_04936_),
    .X(_02594_));
 sky130_fd_sc_hd__nor2_1 _27428_ (.A(net342),
    .B(_04928_),
    .Y(_04937_));
 sky130_vsdinv _27429_ (.A(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_1 _27430_ (.A(_04928_),
    .B(_19666_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _27431_ (.A(_04938_),
    .B(_04939_),
    .Y(_02355_));
 sky130_vsdinv _27432_ (.A(_02356_),
    .Y(_04940_));
 sky130_fd_sc_hd__nor2_2 _27433_ (.A(_20431_),
    .B(_04940_),
    .Y(_04941_));
 sky130_vsdinv _27434_ (.A(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _27435_ (.A(_20431_),
    .B(_04940_),
    .Y(_04943_));
 sky130_fd_sc_hd__nand2_1 _27436_ (.A(_04942_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__a21oi_2 _27437_ (.A1(_04936_),
    .A2(_04930_),
    .B1(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__and3_1 _27438_ (.A(_04936_),
    .B(_04930_),
    .C(_04944_),
    .X(_04946_));
 sky130_fd_sc_hd__nor2_1 _27439_ (.A(_04945_),
    .B(_04946_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_1 _27440_ (.A(_04938_),
    .B(net343),
    .Y(_04947_));
 sky130_fd_sc_hd__nand2_1 _27441_ (.A(_04937_),
    .B(_02357_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _27442_ (.A(_04947_),
    .B(_04948_),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_1 _27443_ (.A(_20051_),
    .B(_02359_),
    .Y(_04949_));
 sky130_fd_sc_hd__nand2_1 _27444_ (.A(_20051_),
    .B(_02359_),
    .Y(_04950_));
 sky130_vsdinv _27445_ (.A(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__nor2_2 _27446_ (.A(_04949_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__a21oi_1 _27447_ (.A1(_04934_),
    .A2(_04932_),
    .B1(_04931_),
    .Y(_04953_));
 sky130_fd_sc_hd__o21ai_1 _27448_ (.A1(_04944_),
    .A2(_04953_),
    .B1(_04942_),
    .Y(_04954_));
 sky130_fd_sc_hd__or2_1 _27449_ (.A(_04952_),
    .B(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__o21ai_2 _27450_ (.A1(_04941_),
    .A2(_04945_),
    .B1(_04952_),
    .Y(_04956_));
 sky130_fd_sc_hd__and2_1 _27451_ (.A(_04955_),
    .B(_04956_),
    .X(_02596_));
 sky130_fd_sc_hd__nor2_2 _27452_ (.A(net344),
    .B(_04948_),
    .Y(_04957_));
 sky130_fd_sc_hd__and2_1 _27453_ (.A(_04948_),
    .B(_19664_),
    .X(_04958_));
 sky130_fd_sc_hd__or2_1 _27454_ (.A(_04957_),
    .B(_04958_),
    .X(_02361_));
 sky130_vsdinv _27455_ (.A(_02362_),
    .Y(_04959_));
 sky130_fd_sc_hd__nor2_2 _27456_ (.A(_20445_),
    .B(_04959_),
    .Y(_04960_));
 sky130_vsdinv _27457_ (.A(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand2_1 _27458_ (.A(_20445_),
    .B(_04959_),
    .Y(_04962_));
 sky130_fd_sc_hd__nand2_2 _27459_ (.A(_04961_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__a21oi_2 _27460_ (.A1(_04956_),
    .A2(_04950_),
    .B1(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__and3_1 _27461_ (.A(_04956_),
    .B(_04950_),
    .C(_04963_),
    .X(_04965_));
 sky130_fd_sc_hd__nor2_1 _27462_ (.A(_04964_),
    .B(_04965_),
    .Y(_02597_));
 sky130_fd_sc_hd__or2_1 _27463_ (.A(_02363_),
    .B(_04957_),
    .X(_04966_));
 sky130_fd_sc_hd__nand2_1 _27464_ (.A(_04957_),
    .B(_02363_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand2_1 _27465_ (.A(_04966_),
    .B(_04967_),
    .Y(_02364_));
 sky130_vsdinv _27466_ (.A(_02365_),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _27467_ (.A(_20776_),
    .B(_04968_),
    .Y(_04969_));
 sky130_vsdinv _27468_ (.A(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2_1 _27469_ (.A(_20776_),
    .B(_04968_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_1 _27470_ (.A(_04970_),
    .B(_04971_),
    .Y(_04972_));
 sky130_vsdinv _27471_ (.A(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__a21oi_2 _27472_ (.A1(_04954_),
    .A2(_04952_),
    .B1(_04951_),
    .Y(_04974_));
 sky130_fd_sc_hd__o21ai_2 _27473_ (.A1(_04963_),
    .A2(_04974_),
    .B1(_04961_),
    .Y(_04975_));
 sky130_fd_sc_hd__nor2_1 _27474_ (.A(_04973_),
    .B(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__and2_1 _27475_ (.A(_04975_),
    .B(_04973_),
    .X(_04977_));
 sky130_fd_sc_hd__nor2_1 _27476_ (.A(_04976_),
    .B(_04977_),
    .Y(_02598_));
 sky130_fd_sc_hd__or2_2 _27477_ (.A(net346),
    .B(_04967_),
    .X(_04978_));
 sky130_fd_sc_hd__nand2_1 _27478_ (.A(_04967_),
    .B(_19663_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _27479_ (.A(_04978_),
    .B(_04979_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _27480_ (.A(net314),
    .B(_02368_),
    .Y(_04980_));
 sky130_vsdinv _27481_ (.A(_02368_),
    .Y(_04981_));
 sky130_fd_sc_hd__nor2_1 _27482_ (.A(_20396_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_2 _27483_ (.A(_04980_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__nor2_1 _27484_ (.A(_04969_),
    .B(_04977_),
    .Y(_04984_));
 sky130_fd_sc_hd__xnor2_1 _27485_ (.A(_04983_),
    .B(_04984_),
    .Y(_02599_));
 sky130_fd_sc_hd__nor2_1 _27486_ (.A(net347),
    .B(_04978_),
    .Y(_04985_));
 sky130_vsdinv _27487_ (.A(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _27488_ (.A(_04978_),
    .B(_19662_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _27489_ (.A(_04986_),
    .B(_04987_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_1 _27490_ (.A(_04973_),
    .B(_04983_),
    .Y(_04988_));
 sky130_fd_sc_hd__o21bai_1 _27491_ (.A1(_04960_),
    .A2(_04964_),
    .B1_N(_04988_),
    .Y(_04989_));
 sky130_vsdinv _27492_ (.A(_04982_),
    .Y(_04990_));
 sky130_fd_sc_hd__o21a_1 _27493_ (.A1(_04980_),
    .A2(_04970_),
    .B1(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _27494_ (.A(_20049_),
    .B(_02371_),
    .Y(_04992_));
 sky130_fd_sc_hd__and2_1 _27495_ (.A(net315),
    .B(_02371_),
    .X(_04993_));
 sky130_fd_sc_hd__nor2_1 _27496_ (.A(_04992_),
    .B(_04993_),
    .Y(_04994_));
 sky130_vsdinv _27497_ (.A(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__a21oi_1 _27498_ (.A1(_04989_),
    .A2(_04991_),
    .B1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__and3_1 _27499_ (.A(_04989_),
    .B(_04995_),
    .C(_04991_),
    .X(_04997_));
 sky130_fd_sc_hd__nor2_1 _27500_ (.A(_04996_),
    .B(_04997_),
    .Y(_02600_));
 sky130_fd_sc_hd__nor2_1 _27501_ (.A(_02372_),
    .B(_04985_),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_1 _27502_ (.A(net348),
    .B(_04986_),
    .Y(_04999_));
 sky130_fd_sc_hd__or2_1 _27503_ (.A(_04998_),
    .B(_04999_),
    .X(_02373_));
 sky130_fd_sc_hd__nor2_1 _27504_ (.A(_20047_),
    .B(_02374_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _27505_ (.A(net316),
    .B(_02374_),
    .Y(_05001_));
 sky130_vsdinv _27506_ (.A(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__nor2_1 _27507_ (.A(_05000_),
    .B(_05002_),
    .Y(_05003_));
 sky130_vsdinv _27508_ (.A(_04991_),
    .Y(_05004_));
 sky130_fd_sc_hd__a31oi_1 _27509_ (.A1(_04975_),
    .A2(_04973_),
    .A3(_04983_),
    .B1(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__o21bai_1 _27510_ (.A1(_04995_),
    .A2(_05005_),
    .B1_N(_04993_),
    .Y(_05006_));
 sky130_fd_sc_hd__or2_1 _27511_ (.A(_05003_),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__o21ai_1 _27512_ (.A1(_04993_),
    .A2(_04996_),
    .B1(_05003_),
    .Y(_05008_));
 sky130_fd_sc_hd__and2_1 _27513_ (.A(_05007_),
    .B(_05008_),
    .X(_02601_));
 sky130_fd_sc_hd__or2_1 _27514_ (.A(_02375_),
    .B(_04999_),
    .X(_05009_));
 sky130_fd_sc_hd__nand2_1 _27515_ (.A(_04999_),
    .B(_02375_),
    .Y(_05010_));
 sky130_fd_sc_hd__nand2_1 _27516_ (.A(_05009_),
    .B(_05010_),
    .Y(_02376_));
 sky130_fd_sc_hd__or2_1 _27517_ (.A(_20046_),
    .B(_02377_),
    .X(_05011_));
 sky130_fd_sc_hd__nand2_1 _27518_ (.A(_20046_),
    .B(_02377_),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_1 _27519_ (.A(_05011_),
    .B(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__a21oi_1 _27520_ (.A1(_05008_),
    .A2(_05001_),
    .B1(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__and3_1 _27521_ (.A(_05008_),
    .B(_05001_),
    .C(_05013_),
    .X(_05015_));
 sky130_fd_sc_hd__nor2_1 _27522_ (.A(_05014_),
    .B(_05015_),
    .Y(_02603_));
 sky130_fd_sc_hd__nor2_1 _27523_ (.A(net351),
    .B(_05010_),
    .Y(_05016_));
 sky130_vsdinv _27524_ (.A(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _27525_ (.A(_05010_),
    .B(_19660_),
    .Y(_05018_));
 sky130_fd_sc_hd__nand2_1 _27526_ (.A(_05017_),
    .B(_05018_),
    .Y(_02379_));
 sky130_fd_sc_hd__nor2_1 _27527_ (.A(_20045_),
    .B(_02380_),
    .Y(_05019_));
 sky130_fd_sc_hd__nand2_1 _27528_ (.A(net319),
    .B(_02380_),
    .Y(_05020_));
 sky130_vsdinv _27529_ (.A(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__nor2_1 _27530_ (.A(_05019_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__a21oi_1 _27531_ (.A1(_05006_),
    .A2(_05003_),
    .B1(_05002_),
    .Y(_05023_));
 sky130_fd_sc_hd__o21ai_1 _27532_ (.A1(_05013_),
    .A2(_05023_),
    .B1(_05012_),
    .Y(_05024_));
 sky130_fd_sc_hd__or2_1 _27533_ (.A(_05022_),
    .B(_05024_),
    .X(_05025_));
 sky130_vsdinv _27534_ (.A(_05012_),
    .Y(_05026_));
 sky130_vsdinv _27535_ (.A(_05022_),
    .Y(_05027_));
 sky130_fd_sc_hd__o21bai_1 _27536_ (.A1(_05026_),
    .A2(_05014_),
    .B1_N(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__and2_1 _27537_ (.A(_05025_),
    .B(_05028_),
    .X(_02604_));
 sky130_fd_sc_hd__nand2_1 _27538_ (.A(_05017_),
    .B(net352),
    .Y(_05029_));
 sky130_fd_sc_hd__nand2_1 _27539_ (.A(_05016_),
    .B(_02381_),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _27540_ (.A(_05029_),
    .B(_05030_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor2_1 _27541_ (.A(_20044_),
    .B(_02383_),
    .Y(_05031_));
 sky130_fd_sc_hd__and2_1 _27542_ (.A(net320),
    .B(_02383_),
    .X(_05032_));
 sky130_fd_sc_hd__or2_1 _27543_ (.A(_05031_),
    .B(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__a21oi_1 _27544_ (.A1(_05028_),
    .A2(_05020_),
    .B1(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__and3_1 _27545_ (.A(_05028_),
    .B(_05020_),
    .C(_05033_),
    .X(_05035_));
 sky130_fd_sc_hd__nor2_1 _27546_ (.A(_05034_),
    .B(_05035_),
    .Y(_02605_));
 sky130_fd_sc_hd__nor2_1 _27547_ (.A(net353),
    .B(_05030_),
    .Y(_05036_));
 sky130_vsdinv _27548_ (.A(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _27549_ (.A(_05030_),
    .B(net353),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _27550_ (.A(_05037_),
    .B(_05038_),
    .Y(_02385_));
 sky130_fd_sc_hd__nor2_2 _27551_ (.A(_20043_),
    .B(_02386_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _27552_ (.A(net321),
    .B(_02386_),
    .Y(_05040_));
 sky130_vsdinv _27553_ (.A(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__nor2_4 _27554_ (.A(_05039_),
    .B(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__a21oi_1 _27555_ (.A1(_05024_),
    .A2(_05022_),
    .B1(_05021_),
    .Y(_05043_));
 sky130_fd_sc_hd__o21bai_2 _27556_ (.A1(_05033_),
    .A2(_05043_),
    .B1_N(_05032_),
    .Y(_05044_));
 sky130_fd_sc_hd__or2_1 _27557_ (.A(_05042_),
    .B(_05044_),
    .X(_05045_));
 sky130_vsdinv _27558_ (.A(_05042_),
    .Y(_05046_));
 sky130_fd_sc_hd__o21bai_1 _27559_ (.A1(_05032_),
    .A2(_05034_),
    .B1_N(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__and2_1 _27560_ (.A(_05045_),
    .B(_05047_),
    .X(_02606_));
 sky130_fd_sc_hd__nand2_1 _27561_ (.A(_05037_),
    .B(net354),
    .Y(_05048_));
 sky130_fd_sc_hd__nand2_1 _27562_ (.A(_05036_),
    .B(_02387_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2_1 _27563_ (.A(_05048_),
    .B(_05049_),
    .Y(_02388_));
 sky130_fd_sc_hd__or2_1 _27564_ (.A(net322),
    .B(_02389_),
    .X(_05050_));
 sky130_fd_sc_hd__nand2_1 _27565_ (.A(net322),
    .B(_02389_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand2_1 _27566_ (.A(_05050_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__a21oi_4 _27567_ (.A1(_05044_),
    .A2(_05042_),
    .B1(_05041_),
    .Y(_05053_));
 sky130_fd_sc_hd__or2_1 _27568_ (.A(_05052_),
    .B(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__nand2_1 _27569_ (.A(_05053_),
    .B(_05052_),
    .Y(_05055_));
 sky130_fd_sc_hd__and2_1 _27570_ (.A(_05054_),
    .B(_05055_),
    .X(_02607_));
 sky130_fd_sc_hd__or2_1 _27571_ (.A(_19659_),
    .B(_05049_),
    .X(_05056_));
 sky130_fd_sc_hd__nand2_1 _27572_ (.A(_05049_),
    .B(_19659_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand2_1 _27573_ (.A(_05056_),
    .B(_05057_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_2 _27574_ (.A(_20040_),
    .B(_02392_),
    .Y(_05058_));
 sky130_fd_sc_hd__and2_1 _27575_ (.A(_20040_),
    .B(_02392_),
    .X(_05059_));
 sky130_fd_sc_hd__nor2_1 _27576_ (.A(_05058_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _27577_ (.A(_05054_),
    .B(_05051_),
    .Y(_05061_));
 sky130_fd_sc_hd__xor2_1 _27578_ (.A(_05060_),
    .B(_05061_),
    .X(_02608_));
 sky130_fd_sc_hd__or2_1 _27579_ (.A(_19657_),
    .B(_05056_),
    .X(_05062_));
 sky130_fd_sc_hd__nand2_1 _27580_ (.A(_05056_),
    .B(_19657_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _27581_ (.A(_05062_),
    .B(_05063_),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_1 _27582_ (.A(_20039_),
    .B(_02395_),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_1 _27583_ (.A(_20039_),
    .B(_02395_),
    .Y(_05065_));
 sky130_fd_sc_hd__nand2_1 _27584_ (.A(_05064_),
    .B(_05065_),
    .Y(_05066_));
 sky130_vsdinv _27585_ (.A(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__or3_4 _27586_ (.A(_05058_),
    .B(_05059_),
    .C(_05052_),
    .X(_05068_));
 sky130_fd_sc_hd__o21bai_1 _27587_ (.A1(_05051_),
    .A2(_05058_),
    .B1_N(_05059_),
    .Y(_05069_));
 sky130_fd_sc_hd__o21bai_4 _27588_ (.A1(_05068_),
    .A2(_05053_),
    .B1_N(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__or2_1 _27589_ (.A(_05067_),
    .B(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__nand2_1 _27590_ (.A(_05070_),
    .B(_05067_),
    .Y(_05072_));
 sky130_fd_sc_hd__and2_1 _27591_ (.A(_05071_),
    .B(_05072_),
    .X(_02609_));
 sky130_fd_sc_hd__nor2_1 _27592_ (.A(_19656_),
    .B(_05062_),
    .Y(_05073_));
 sky130_vsdinv _27593_ (.A(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand2_1 _27594_ (.A(_05062_),
    .B(_19656_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand2_1 _27595_ (.A(_05074_),
    .B(_05075_),
    .Y(_02397_));
 sky130_fd_sc_hd__nor2_1 _27596_ (.A(net325),
    .B(_02398_),
    .Y(_05076_));
 sky130_vsdinv _27597_ (.A(_02398_),
    .Y(_05077_));
 sky130_fd_sc_hd__nor2_1 _27598_ (.A(_20522_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__nor2_2 _27599_ (.A(_05076_),
    .B(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_1 _27600_ (.A(_05072_),
    .B(_05065_),
    .Y(_05080_));
 sky130_fd_sc_hd__xor2_1 _27601_ (.A(_05079_),
    .B(_05080_),
    .X(_02610_));
 sky130_fd_sc_hd__nand2_1 _27602_ (.A(_05074_),
    .B(net358),
    .Y(_05081_));
 sky130_fd_sc_hd__nand2_1 _27603_ (.A(_05073_),
    .B(_02399_),
    .Y(_05082_));
 sky130_fd_sc_hd__nand2_1 _27604_ (.A(_05081_),
    .B(_05082_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _27605_ (.A(_20038_),
    .B(_02401_),
    .Y(_05083_));
 sky130_vsdinv _27606_ (.A(_02401_),
    .Y(_05084_));
 sky130_fd_sc_hd__nor2_2 _27607_ (.A(_20505_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__or2_1 _27608_ (.A(_05083_),
    .B(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__nand2_1 _27609_ (.A(_05067_),
    .B(_05079_),
    .Y(_05087_));
 sky130_vsdinv _27610_ (.A(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__o21ba_1 _27611_ (.A1(_05065_),
    .A2(_05076_),
    .B1_N(_05078_),
    .X(_05089_));
 sky130_fd_sc_hd__a21boi_4 _27612_ (.A1(_05070_),
    .A2(_05088_),
    .B1_N(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__xor2_1 _27613_ (.A(_05086_),
    .B(_05090_),
    .X(_02611_));
 sky130_fd_sc_hd__nor2_1 _27614_ (.A(_19655_),
    .B(_05082_),
    .Y(_05091_));
 sky130_vsdinv _27615_ (.A(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand2_1 _27616_ (.A(_05082_),
    .B(_19655_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _27617_ (.A(_05092_),
    .B(_05093_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _27618_ (.A(_20037_),
    .B(_02404_),
    .Y(_05094_));
 sky130_vsdinv _27619_ (.A(_02404_),
    .Y(_05095_));
 sky130_fd_sc_hd__nor2_2 _27620_ (.A(_20518_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__nor2_1 _27621_ (.A(_05094_),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__o21bai_2 _27622_ (.A1(_05083_),
    .A2(_05090_),
    .B1_N(_05085_),
    .Y(_05098_));
 sky130_fd_sc_hd__xor2_1 _27623_ (.A(_05097_),
    .B(_05098_),
    .X(_02612_));
 sky130_fd_sc_hd__nand2_1 _27624_ (.A(_05092_),
    .B(net361),
    .Y(_05099_));
 sky130_fd_sc_hd__nand2_1 _27625_ (.A(_05091_),
    .B(_02405_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _27626_ (.A(_05099_),
    .B(_05100_),
    .Y(_02406_));
 sky130_vsdinv _27627_ (.A(_05094_),
    .Y(_05101_));
 sky130_fd_sc_hd__a21oi_2 _27628_ (.A1(_05098_),
    .A2(_05101_),
    .B1(_05096_),
    .Y(_05102_));
 sky130_fd_sc_hd__nor2_1 _27629_ (.A(_20036_),
    .B(_02407_),
    .Y(_05103_));
 sky130_vsdinv _27630_ (.A(_02407_),
    .Y(_05104_));
 sky130_fd_sc_hd__nor2_2 _27631_ (.A(_20529_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__nor2_1 _27632_ (.A(_05103_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2_1 _27633_ (.A(_05102_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__a21oi_2 _27634_ (.A1(_05047_),
    .A2(_05040_),
    .B1(_05068_),
    .Y(_05108_));
 sky130_fd_sc_hd__o21bai_2 _27635_ (.A1(_05069_),
    .A2(_05108_),
    .B1_N(_05087_),
    .Y(_05109_));
 sky130_fd_sc_hd__a22oi_2 _27636_ (.A1(_20505_),
    .A2(_05084_),
    .B1(_05109_),
    .B2(_05089_),
    .Y(_05110_));
 sky130_fd_sc_hd__o22ai_2 _27637_ (.A1(_20037_),
    .A2(_02404_),
    .B1(_05085_),
    .B2(_05110_),
    .Y(_05111_));
 sky130_vsdinv _27638_ (.A(_05096_),
    .Y(_05112_));
 sky130_fd_sc_hd__a21o_1 _27639_ (.A1(_05111_),
    .A2(_05112_),
    .B1(_05106_),
    .X(_05113_));
 sky130_fd_sc_hd__nand2_1 _27640_ (.A(_05107_),
    .B(_05113_),
    .Y(_02614_));
 sky130_fd_sc_hd__xor2_1 _27641_ (.A(net362),
    .B(_05100_),
    .X(_02408_));
 sky130_fd_sc_hd__nor2_1 _27642_ (.A(_02409_),
    .B(_18667_),
    .Y(_05114_));
 sky130_fd_sc_hd__and2_1 _27643_ (.A(_18667_),
    .B(_02409_),
    .X(_05115_));
 sky130_fd_sc_hd__a22oi_1 _27644_ (.A1(_20529_),
    .A2(_05104_),
    .B1(_05111_),
    .B2(_05112_),
    .Y(_05116_));
 sky130_fd_sc_hd__o22ai_1 _27645_ (.A1(_05114_),
    .A2(_05115_),
    .B1(_05105_),
    .B2(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__or3_2 _27646_ (.A(_05114_),
    .B(_05105_),
    .C(_05115_),
    .X(_05118_));
 sky130_fd_sc_hd__o21bai_1 _27647_ (.A1(_05103_),
    .A2(_05102_),
    .B1_N(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__nand2_1 _27648_ (.A(_05117_),
    .B(_05119_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _27649_ (.A(_19939_),
    .B(_20175_),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _27650_ (.A(_19935_),
    .B(_20178_),
    .Y(_05121_));
 sky130_fd_sc_hd__nor2_4 _27651_ (.A(_05120_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__and2_2 _27652_ (.A(_05120_),
    .B(_05121_),
    .X(_05123_));
 sky130_fd_sc_hd__nor2_8 _27653_ (.A(_05122_),
    .B(_05123_),
    .Y(_02624_));
 sky130_vsdinv _27654_ (.A(_05122_),
    .Y(_05124_));
 sky130_fd_sc_hd__buf_6 _27655_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05125_));
 sky130_fd_sc_hd__clkinv_8 _27656_ (.A(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__clkbuf_4 _27657_ (.A(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__nor2_2 _27658_ (.A(net470),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__nand2_4 _27659_ (.A(_19930_),
    .B(_19933_),
    .Y(_05129_));
 sky130_fd_sc_hd__buf_6 _27660_ (.A(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__buf_4 _27661_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05131_));
 sky130_vsdinv _27662_ (.A(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__or2_1 _27663_ (.A(_05130_),
    .B(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__a22o_1 _27664_ (.A1(_19932_),
    .A2(_20178_),
    .B1(_19935_),
    .B2(_20175_),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_2 _27665_ (.A1(_04841_),
    .A2(_05133_),
    .B1(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__xor2_2 _27666_ (.A(_05128_),
    .B(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__nor2_2 _27667_ (.A(_05124_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__and2_1 _27668_ (.A(_05136_),
    .B(_05124_),
    .X(_05138_));
 sky130_fd_sc_hd__nor2_1 _27669_ (.A(_05137_),
    .B(_05138_),
    .Y(_02625_));
 sky130_fd_sc_hd__buf_6 _27670_ (.A(_19930_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_4 _27671_ (.A(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__buf_6 _27672_ (.A(_19933_),
    .X(_05141_));
 sky130_fd_sc_hd__buf_4 _27673_ (.A(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__buf_4 _27674_ (.A(_05125_),
    .X(_05143_));
 sky130_fd_sc_hd__buf_6 _27675_ (.A(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__buf_6 _27676_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05145_));
 sky130_fd_sc_hd__buf_6 _27677_ (.A(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__buf_6 _27678_ (.A(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__and4_2 _27679_ (.A(_05140_),
    .B(_05142_),
    .C(_05144_),
    .D(_05147_),
    .X(_05148_));
 sky130_vsdinv _27680_ (.A(_05140_),
    .Y(_05149_));
 sky130_vsdinv _27681_ (.A(_19933_),
    .Y(_05150_));
 sky130_fd_sc_hd__buf_6 _27682_ (.A(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__o22a_1 _27683_ (.A1(_05149_),
    .A2(_05132_),
    .B1(_05151_),
    .B2(_05127_),
    .X(_05152_));
 sky130_vsdinv _27684_ (.A(\pcpi_mul.rs2[3] ),
    .Y(_05153_));
 sky130_fd_sc_hd__buf_6 _27685_ (.A(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_4 _27686_ (.A(_05154_),
    .B(_04839_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21bai_2 _27687_ (.A1(_05148_),
    .A2(_05152_),
    .B1_N(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__a22o_2 _27688_ (.A1(_19932_),
    .A2(_20175_),
    .B1(_19935_),
    .B2(_20172_),
    .X(_05157_));
 sky130_fd_sc_hd__nand3b_4 _27689_ (.A_N(_05148_),
    .B(_05157_),
    .C(_05155_),
    .Y(_05158_));
 sky130_fd_sc_hd__nand2_1 _27690_ (.A(_05156_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_2 _27691_ (.A(_19939_),
    .B(_20169_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_2 _27692_ (.A(_05159_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand3b_4 _27693_ (.A_N(_05160_),
    .B(_05156_),
    .C(_05158_),
    .Y(_05162_));
 sky130_fd_sc_hd__a2bb2o_2 _27694_ (.A1_N(_04840_),
    .A2_N(_05133_),
    .B1(_05128_),
    .B2(_05134_),
    .X(_05163_));
 sky130_fd_sc_hd__a21o_1 _27695_ (.A1(_05161_),
    .A2(_05162_),
    .B1(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__nand3_1 _27696_ (.A(_05161_),
    .B(_05162_),
    .C(_05163_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_1 _27697_ (.A(_05164_),
    .B(_05165_),
    .Y(_05166_));
 sky130_vsdinv _27698_ (.A(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__nor2_1 _27699_ (.A(_05137_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_1 _27700_ (.A(_05167_),
    .B(_05137_),
    .Y(_05169_));
 sky130_vsdinv _27701_ (.A(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__nor2_1 _27702_ (.A(_05168_),
    .B(_05170_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand2_1 _27703_ (.A(_05169_),
    .B(_05165_),
    .Y(_05171_));
 sky130_fd_sc_hd__a21oi_4 _27704_ (.A1(_05155_),
    .A2(_05157_),
    .B1(_05148_),
    .Y(_05172_));
 sky130_fd_sc_hd__buf_4 _27705_ (.A(_19930_),
    .X(_05173_));
 sky130_fd_sc_hd__buf_4 _27706_ (.A(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__buf_6 _27707_ (.A(_05141_),
    .X(_05175_));
 sky130_fd_sc_hd__buf_6 _27708_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_4 _27709_ (.A(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__buf_4 _27710_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05178_));
 sky130_fd_sc_hd__buf_6 _27711_ (.A(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__and4_2 _27712_ (.A(_05174_),
    .B(_05175_),
    .C(_05177_),
    .D(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_4 _27713_ (.A(_05143_),
    .X(_05181_));
 sky130_fd_sc_hd__buf_6 _27714_ (.A(_20167_),
    .X(_05182_));
 sky130_fd_sc_hd__buf_4 _27715_ (.A(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__a22o_1 _27716_ (.A1(_05174_),
    .A2(_05181_),
    .B1(_05142_),
    .B2(_05183_),
    .X(_05184_));
 sky130_vsdinv _27717_ (.A(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__buf_6 _27718_ (.A(_05153_),
    .X(_05186_));
 sky130_fd_sc_hd__nor2_2 _27719_ (.A(_05186_),
    .B(_05132_),
    .Y(_05187_));
 sky130_fd_sc_hd__o21bai_2 _27720_ (.A1(_05180_),
    .A2(_05185_),
    .B1_N(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand3b_4 _27721_ (.A_N(_05180_),
    .B(_05184_),
    .C(_05187_),
    .Y(_05189_));
 sky130_fd_sc_hd__nand2_1 _27722_ (.A(_05188_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand2_1 _27723_ (.A(_19925_),
    .B(_20177_),
    .Y(_05191_));
 sky130_fd_sc_hd__clkbuf_8 _27724_ (.A(_19936_),
    .X(_05192_));
 sky130_fd_sc_hd__nand2_1 _27725_ (.A(_05192_),
    .B(_20165_),
    .Y(_05193_));
 sky130_fd_sc_hd__nor2_2 _27726_ (.A(_05191_),
    .B(_05193_),
    .Y(_05194_));
 sky130_vsdinv _27727_ (.A(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__nand2_1 _27728_ (.A(_05191_),
    .B(_05193_),
    .Y(_05196_));
 sky130_fd_sc_hd__nand2_1 _27729_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__nand2_1 _27730_ (.A(_05190_),
    .B(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand3b_4 _27731_ (.A_N(_05197_),
    .B(_05188_),
    .C(_05189_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2_2 _27732_ (.A(_05198_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2_1 _27733_ (.A(_05200_),
    .B(_05162_),
    .Y(_05201_));
 sky130_fd_sc_hd__nor2_1 _27734_ (.A(_05160_),
    .B(_05159_),
    .Y(_05202_));
 sky130_fd_sc_hd__nand3_2 _27735_ (.A(_05202_),
    .B(_05198_),
    .C(_05199_),
    .Y(_05203_));
 sky130_fd_sc_hd__nand2_1 _27736_ (.A(_05201_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__or2_1 _27737_ (.A(_05172_),
    .B(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__nand2_1 _27738_ (.A(_05204_),
    .B(_05172_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _27739_ (.A(_05205_),
    .B(_05206_),
    .Y(_05207_));
 sky130_vsdinv _27740_ (.A(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__or2_1 _27741_ (.A(_05171_),
    .B(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__nand2_1 _27742_ (.A(_05208_),
    .B(_05171_),
    .Y(_05210_));
 sky130_fd_sc_hd__and2_1 _27743_ (.A(_05209_),
    .B(_05210_),
    .X(_02627_));
 sky130_fd_sc_hd__buf_6 _27744_ (.A(_19923_),
    .X(_05211_));
 sky130_fd_sc_hd__nand2_4 _27745_ (.A(_05211_),
    .B(_05131_),
    .Y(_05212_));
 sky130_fd_sc_hd__buf_8 _27746_ (.A(_19919_),
    .X(_05213_));
 sky130_fd_sc_hd__buf_4 _27747_ (.A(_20176_),
    .X(_05214_));
 sky130_fd_sc_hd__nand2_4 _27748_ (.A(_05213_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__nor2_8 _27749_ (.A(_05212_),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__clkbuf_2 _27750_ (.A(_19936_),
    .X(_05217_));
 sky130_fd_sc_hd__buf_4 _27751_ (.A(_20161_),
    .X(_05218_));
 sky130_fd_sc_hd__nand2_2 _27752_ (.A(net469),
    .B(_05218_),
    .Y(_05219_));
 sky130_vsdinv _27753_ (.A(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand2_2 _27754_ (.A(_05212_),
    .B(_05215_),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_1 _27755_ (.A(_05220_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__a22oi_4 _27756_ (.A1(_19920_),
    .A2(_20177_),
    .B1(_19925_),
    .B2(_05146_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ai_2 _27757_ (.A1(_05223_),
    .A2(_05216_),
    .B1(_05219_),
    .Y(_05224_));
 sky130_fd_sc_hd__o211ai_4 _27758_ (.A1(_05216_),
    .A2(_05222_),
    .B1(_05194_),
    .C1(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__o21ai_2 _27759_ (.A1(_05223_),
    .A2(_05216_),
    .B1(_05220_),
    .Y(_05226_));
 sky130_fd_sc_hd__clkbuf_4 _27760_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05227_));
 sky130_fd_sc_hd__buf_6 _27761_ (.A(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__clkbuf_8 _27762_ (.A(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__buf_6 _27763_ (.A(_04838_),
    .X(_05230_));
 sky130_fd_sc_hd__nand3b_2 _27764_ (.A_N(_05212_),
    .B(_05229_),
    .C(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand3_2 _27765_ (.A(_05231_),
    .B(_05221_),
    .C(_05219_),
    .Y(_05232_));
 sky130_fd_sc_hd__nand3_4 _27766_ (.A(_05226_),
    .B(_05232_),
    .C(_05195_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_1 _27767_ (.A(_05225_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__buf_4 _27768_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05235_));
 sky130_fd_sc_hd__buf_6 _27769_ (.A(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_4 _27770_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05237_));
 sky130_fd_sc_hd__buf_6 _27771_ (.A(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__a22oi_4 _27772_ (.A1(_05236_),
    .A2(_05177_),
    .B1(_05175_),
    .B2(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__clkbuf_4 _27773_ (.A(_19930_),
    .X(_05240_));
 sky130_fd_sc_hd__buf_2 _27774_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05241_));
 sky130_fd_sc_hd__buf_4 _27775_ (.A(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__buf_4 _27776_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05243_));
 sky130_fd_sc_hd__buf_6 _27777_ (.A(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__buf_6 _27778_ (.A(_20167_),
    .X(_05245_));
 sky130_fd_sc_hd__and4_4 _27779_ (.A(_05240_),
    .B(_05242_),
    .C(_05244_),
    .D(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__buf_6 _27780_ (.A(_19927_),
    .X(_05247_));
 sky130_fd_sc_hd__nand2_4 _27781_ (.A(_05247_),
    .B(_20171_),
    .Y(_05248_));
 sky130_fd_sc_hd__o21bai_1 _27782_ (.A1(_05239_),
    .A2(_05246_),
    .B1_N(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__buf_6 _27783_ (.A(_05150_),
    .X(_05250_));
 sky130_fd_sc_hd__buf_6 _27784_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05251_));
 sky130_vsdinv _27785_ (.A(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__buf_6 _27786_ (.A(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__nand2_2 _27787_ (.A(_05173_),
    .B(_05182_),
    .Y(_05254_));
 sky130_fd_sc_hd__o21ai_4 _27788_ (.A1(_05250_),
    .A2(_05253_),
    .B1(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__nand3b_4 _27789_ (.A_N(_05254_),
    .B(_05175_),
    .C(_05238_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand3_2 _27790_ (.A(_05255_),
    .B(_05256_),
    .C(_05248_),
    .Y(_05257_));
 sky130_fd_sc_hd__and2_1 _27791_ (.A(_05249_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__nand2_1 _27792_ (.A(_05234_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__nand2_2 _27793_ (.A(_05249_),
    .B(_05257_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand3_2 _27794_ (.A(_05225_),
    .B(_05233_),
    .C(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__nand3b_4 _27795_ (.A_N(_05199_),
    .B(_05259_),
    .C(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2_1 _27796_ (.A(_05234_),
    .B(_05260_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand3_2 _27797_ (.A(_05258_),
    .B(_05225_),
    .C(_05233_),
    .Y(_05264_));
 sky130_fd_sc_hd__nand3_4 _27798_ (.A(_05263_),
    .B(_05264_),
    .C(_05199_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_1 _27799_ (.A(_05262_),
    .B(_05265_),
    .Y(_05266_));
 sky130_vsdinv _27800_ (.A(_05189_),
    .Y(_05267_));
 sky130_fd_sc_hd__nor2_4 _27801_ (.A(_05180_),
    .B(_05267_),
    .Y(_05268_));
 sky130_vsdinv _27802_ (.A(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__nand2_2 _27803_ (.A(_05266_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand3_4 _27804_ (.A(_05262_),
    .B(_05265_),
    .C(_05268_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_1 _27805_ (.A(_05203_),
    .B(_05172_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2_2 _27806_ (.A(_05272_),
    .B(_05201_),
    .Y(_05273_));
 sky130_fd_sc_hd__a21oi_4 _27807_ (.A1(_05270_),
    .A2(_05271_),
    .B1(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__o2111ai_4 _27808_ (.A1(_05172_),
    .A2(_05200_),
    .B1(_05162_),
    .C1(_05161_),
    .D1(_05163_),
    .Y(_05275_));
 sky130_fd_sc_hd__a21oi_1 _27809_ (.A1(_05172_),
    .A2(_05204_),
    .B1(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand3_2 _27810_ (.A(_05270_),
    .B(_05273_),
    .C(_05271_),
    .Y(_05277_));
 sky130_fd_sc_hd__and2_1 _27811_ (.A(_05276_),
    .B(_05277_),
    .X(_05278_));
 sky130_vsdinv _27812_ (.A(_19918_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_2 _27813_ (.A(_05256_),
    .B(_05248_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_4 _27814_ (.A(_19927_),
    .B(_05245_),
    .Y(_05281_));
 sky130_fd_sc_hd__buf_6 _27815_ (.A(_19930_),
    .X(_05282_));
 sky130_fd_sc_hd__clkbuf_8 _27816_ (.A(_05251_),
    .X(_05283_));
 sky130_fd_sc_hd__buf_6 _27817_ (.A(_19933_),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_8 _27818_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05285_));
 sky130_fd_sc_hd__buf_6 _27819_ (.A(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__a22oi_4 _27820_ (.A1(_05282_),
    .A2(_05283_),
    .B1(_05284_),
    .B2(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__clkbuf_4 _27821_ (.A(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__buf_6 _27822_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05289_));
 sky130_fd_sc_hd__and4_1 _27823_ (.A(_05235_),
    .B(_05241_),
    .C(_05289_),
    .D(_05237_),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_4 _27824_ (.A(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__nor3_4 _27825_ (.A(_05281_),
    .B(_05288_),
    .C(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__o21a_1 _27826_ (.A1(_05288_),
    .A2(_05291_),
    .B1(_05281_),
    .X(_05293_));
 sky130_fd_sc_hd__buf_4 _27827_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05294_));
 sky130_vsdinv _27828_ (.A(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__buf_6 _27829_ (.A(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__buf_6 _27830_ (.A(_05145_),
    .X(_05297_));
 sky130_fd_sc_hd__buf_6 _27831_ (.A(_19924_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_4 _27832_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05299_));
 sky130_fd_sc_hd__buf_6 _27833_ (.A(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__a22oi_4 _27834_ (.A1(_05213_),
    .A2(_05297_),
    .B1(_05298_),
    .B2(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__buf_6 _27835_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05302_));
 sky130_fd_sc_hd__nand3_4 _27836_ (.A(_05302_),
    .B(_19924_),
    .C(_05145_),
    .Y(_05303_));
 sky130_fd_sc_hd__nor2_4 _27837_ (.A(_05126_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__o22ai_4 _27838_ (.A1(net470),
    .A2(_05296_),
    .B1(_05301_),
    .B2(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__o21ai_2 _27839_ (.A1(_05219_),
    .A2(_05223_),
    .B1(_05231_),
    .Y(_05306_));
 sky130_fd_sc_hd__buf_4 _27840_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05307_));
 sky130_fd_sc_hd__buf_4 _27841_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05308_));
 sky130_fd_sc_hd__nand2_2 _27842_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 sky130_vsdinv _27843_ (.A(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__buf_6 _27844_ (.A(_05227_),
    .X(_05311_));
 sky130_fd_sc_hd__buf_6 _27845_ (.A(_19923_),
    .X(_05312_));
 sky130_fd_sc_hd__buf_6 _27846_ (.A(_05125_),
    .X(_05313_));
 sky130_fd_sc_hd__a22o_2 _27847_ (.A1(_05311_),
    .A2(_05131_),
    .B1(_05312_),
    .B2(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__o211ai_2 _27848_ (.A1(_05127_),
    .A2(_05303_),
    .B1(_05310_),
    .C1(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand3_4 _27849_ (.A(_05305_),
    .B(_05306_),
    .C(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21ai_2 _27850_ (.A1(_05301_),
    .A2(_05304_),
    .B1(_05310_),
    .Y(_05317_));
 sky130_fd_sc_hd__a21oi_2 _27851_ (.A1(_05220_),
    .A2(_05221_),
    .B1(_05216_),
    .Y(_05318_));
 sky130_fd_sc_hd__o211ai_2 _27852_ (.A1(_05127_),
    .A2(_05303_),
    .B1(_05309_),
    .C1(_05314_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand3_4 _27853_ (.A(_05317_),
    .B(_05318_),
    .C(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__a2bb2oi_2 _27854_ (.A1_N(_05292_),
    .A2_N(_05293_),
    .B1(_05316_),
    .B2(_05320_),
    .Y(_05321_));
 sky130_vsdinv _27855_ (.A(_05281_),
    .Y(_05322_));
 sky130_fd_sc_hd__nor3_1 _27856_ (.A(_05322_),
    .B(_05288_),
    .C(_05291_),
    .Y(_05323_));
 sky130_fd_sc_hd__o21a_1 _27857_ (.A1(_05288_),
    .A2(_05291_),
    .B1(_05322_),
    .X(_05324_));
 sky130_fd_sc_hd__o211a_1 _27858_ (.A1(_05323_),
    .A2(_05324_),
    .B1(_05316_),
    .C1(_05320_),
    .X(_05325_));
 sky130_fd_sc_hd__a21boi_4 _27859_ (.A1(_05260_),
    .A2(_05233_),
    .B1_N(_05225_),
    .Y(_05326_));
 sky130_fd_sc_hd__o21ai_4 _27860_ (.A1(_05321_),
    .A2(_05325_),
    .B1(_05326_),
    .Y(_05327_));
 sky130_vsdinv _27861_ (.A(_05287_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand3b_1 _27862_ (.A_N(_05290_),
    .B(_05328_),
    .C(_05281_),
    .Y(_05329_));
 sky130_fd_sc_hd__o21ai_1 _27863_ (.A1(_05287_),
    .A2(_05291_),
    .B1(_05322_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _27864_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a21o_1 _27865_ (.A1(_05320_),
    .A2(_05316_),
    .B1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__nand2_1 _27866_ (.A(_05233_),
    .B(_05260_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_1 _27867_ (.A(_05333_),
    .B(_05225_),
    .Y(_05334_));
 sky130_fd_sc_hd__nand3_2 _27868_ (.A(_05331_),
    .B(_05320_),
    .C(_05316_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand3_4 _27869_ (.A(_05332_),
    .B(_05334_),
    .C(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__a22oi_4 _27870_ (.A1(_05255_),
    .A2(_05280_),
    .B1(_05327_),
    .B2(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__nor2_4 _27871_ (.A(_05248_),
    .B(_05239_),
    .Y(_05338_));
 sky130_fd_sc_hd__o211a_1 _27872_ (.A1(_05246_),
    .A2(_05338_),
    .B1(_05336_),
    .C1(_05327_),
    .X(_05339_));
 sky130_fd_sc_hd__o22ai_4 _27873_ (.A1(_05279_),
    .A2(_04841_),
    .B1(_05337_),
    .B2(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__nand2_2 _27874_ (.A(_05327_),
    .B(_05336_),
    .Y(_05341_));
 sky130_fd_sc_hd__nor2_8 _27875_ (.A(_05246_),
    .B(_05338_),
    .Y(_05342_));
 sky130_fd_sc_hd__nand2_2 _27876_ (.A(_05341_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__nand3b_4 _27877_ (.A_N(_05342_),
    .B(_05327_),
    .C(_05336_),
    .Y(_05344_));
 sky130_fd_sc_hd__nor2_4 _27878_ (.A(_05279_),
    .B(_04841_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand3_4 _27879_ (.A(_05343_),
    .B(_05344_),
    .C(_05345_),
    .Y(_05346_));
 sky130_vsdinv _27880_ (.A(_05262_),
    .Y(_05347_));
 sky130_fd_sc_hd__and2_1 _27881_ (.A(_05265_),
    .B(_05269_),
    .X(_05348_));
 sky130_fd_sc_hd__or2_2 _27882_ (.A(_05347_),
    .B(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__a21oi_2 _27883_ (.A1(_05340_),
    .A2(_05346_),
    .B1(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__o211a_2 _27884_ (.A1(_05347_),
    .A2(_05348_),
    .B1(_05346_),
    .C1(_05340_),
    .X(_05351_));
 sky130_fd_sc_hd__o22ai_2 _27885_ (.A1(_05274_),
    .A2(_05278_),
    .B1(_05350_),
    .B2(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__a21o_1 _27886_ (.A1(_05340_),
    .A2(_05346_),
    .B1(_05349_),
    .X(_05353_));
 sky130_fd_sc_hd__a21oi_1 _27887_ (.A1(_05276_),
    .A2(_05277_),
    .B1(_05274_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand3_4 _27888_ (.A(_05349_),
    .B(_05340_),
    .C(_05346_),
    .Y(_05355_));
 sky130_fd_sc_hd__nand3_2 _27889_ (.A(_05353_),
    .B(_05354_),
    .C(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__a21o_1 _27890_ (.A1(_05270_),
    .A2(_05271_),
    .B1(_05273_),
    .X(_05357_));
 sky130_fd_sc_hd__nand2_1 _27891_ (.A(_05357_),
    .B(_05277_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand3b_2 _27892_ (.A_N(_05358_),
    .B(_05208_),
    .C(_05170_),
    .Y(_05359_));
 sky130_fd_sc_hd__a21oi_2 _27893_ (.A1(_05352_),
    .A2(_05356_),
    .B1(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__and3_1 _27894_ (.A(_05359_),
    .B(_05352_),
    .C(_05356_),
    .X(_05361_));
 sky130_fd_sc_hd__nor2_1 _27895_ (.A(_05360_),
    .B(_05361_),
    .Y(_02683_));
 sky130_fd_sc_hd__and3_1 _27896_ (.A(_05353_),
    .B(_05355_),
    .C(_05278_),
    .X(_05362_));
 sky130_fd_sc_hd__a21oi_1 _27897_ (.A1(_05353_),
    .A2(_05274_),
    .B1(_05351_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _27898_ (.A(_05331_),
    .B(_05320_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_2 _27899_ (.A(_05364_),
    .B(_05316_),
    .Y(_05365_));
 sky130_fd_sc_hd__buf_6 _27900_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05366_));
 sky130_fd_sc_hd__buf_6 _27901_ (.A(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__a22oi_4 _27902_ (.A1(_05228_),
    .A2(_05313_),
    .B1(_05367_),
    .B2(_05182_),
    .Y(_05368_));
 sky130_fd_sc_hd__clkinv_16 _27903_ (.A(\pcpi_mul.rs1[3] ),
    .Y(_05369_));
 sky130_fd_sc_hd__nand3_4 _27904_ (.A(_19919_),
    .B(_19923_),
    .C(_05125_),
    .Y(_05370_));
 sky130_fd_sc_hd__nor2_8 _27905_ (.A(_05369_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__buf_6 _27906_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05372_));
 sky130_fd_sc_hd__nand2_4 _27907_ (.A(_19936_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__o21ai_2 _27908_ (.A1(_05368_),
    .A2(_05371_),
    .B1(_05373_),
    .Y(_05374_));
 sky130_vsdinv _27909_ (.A(_05373_),
    .Y(_05375_));
 sky130_fd_sc_hd__buf_6 _27910_ (.A(_05227_),
    .X(_05376_));
 sky130_fd_sc_hd__buf_6 _27911_ (.A(_19923_),
    .X(_05377_));
 sky130_fd_sc_hd__a22o_2 _27912_ (.A1(_05376_),
    .A2(_05178_),
    .B1(_05377_),
    .B2(_05176_),
    .X(_05378_));
 sky130_fd_sc_hd__o211ai_4 _27913_ (.A1(_05369_),
    .A2(_05370_),
    .B1(_05375_),
    .C1(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__o22ai_4 _27914_ (.A1(_05127_),
    .A2(_05303_),
    .B1(_05309_),
    .B2(_05301_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand3_4 _27915_ (.A(_05374_),
    .B(_05379_),
    .C(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__o21ai_2 _27916_ (.A1(_05368_),
    .A2(_05371_),
    .B1(_05375_),
    .Y(_05382_));
 sky130_fd_sc_hd__a21oi_2 _27917_ (.A1(_05314_),
    .A2(_05310_),
    .B1(_05304_),
    .Y(_05383_));
 sky130_fd_sc_hd__o211ai_4 _27918_ (.A1(_05369_),
    .A2(_05370_),
    .B1(_05373_),
    .C1(_05378_),
    .Y(_05384_));
 sky130_fd_sc_hd__nand3_4 _27919_ (.A(_05382_),
    .B(_05383_),
    .C(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_4 _27920_ (.A(_05247_),
    .B(_20165_),
    .Y(_05386_));
 sky130_fd_sc_hd__buf_4 _27921_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05387_));
 sky130_fd_sc_hd__buf_6 _27922_ (.A(_20161_),
    .X(_05388_));
 sky130_fd_sc_hd__buf_4 _27923_ (.A(_05294_),
    .X(_05389_));
 sky130_fd_sc_hd__a22oi_4 _27924_ (.A1(_05387_),
    .A2(_05388_),
    .B1(_05141_),
    .B2(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__buf_4 _27925_ (.A(_05294_),
    .X(_05391_));
 sky130_fd_sc_hd__buf_4 _27926_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05392_));
 sky130_fd_sc_hd__and4_4 _27927_ (.A(_05387_),
    .B(_05241_),
    .C(_05391_),
    .D(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__nor3_4 _27928_ (.A(_05386_),
    .B(_05390_),
    .C(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__o21a_1 _27929_ (.A1(_05390_),
    .A2(_05393_),
    .B1(_05386_),
    .X(_05395_));
 sky130_fd_sc_hd__o2bb2ai_2 _27930_ (.A1_N(_05381_),
    .A2_N(_05385_),
    .B1(_05394_),
    .B2(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__nor2_2 _27931_ (.A(_05394_),
    .B(_05395_),
    .Y(_05397_));
 sky130_fd_sc_hd__nand3_2 _27932_ (.A(_05397_),
    .B(_05381_),
    .C(_05385_),
    .Y(_05398_));
 sky130_fd_sc_hd__nand3_4 _27933_ (.A(_05365_),
    .B(_05396_),
    .C(_05398_),
    .Y(_05399_));
 sky130_vsdinv _27934_ (.A(_05320_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21a_1 _27935_ (.A1(_05292_),
    .A2(_05293_),
    .B1(_05316_),
    .X(_05401_));
 sky130_fd_sc_hd__a2bb2oi_2 _27936_ (.A1_N(_05394_),
    .A2_N(_05395_),
    .B1(_05381_),
    .B2(_05385_),
    .Y(_05402_));
 sky130_vsdinv _27937_ (.A(_05386_),
    .Y(_05403_));
 sky130_fd_sc_hd__nor3_1 _27938_ (.A(_05403_),
    .B(_05390_),
    .C(_05393_),
    .Y(_05404_));
 sky130_fd_sc_hd__o21a_1 _27939_ (.A1(_05390_),
    .A2(_05393_),
    .B1(_05403_),
    .X(_05405_));
 sky130_fd_sc_hd__o211a_1 _27940_ (.A1(_05404_),
    .A2(_05405_),
    .B1(_05381_),
    .C1(_05385_),
    .X(_05406_));
 sky130_fd_sc_hd__o22ai_4 _27941_ (.A1(_05400_),
    .A2(_05401_),
    .B1(_05402_),
    .B2(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__nor2_4 _27942_ (.A(_05322_),
    .B(_05291_),
    .Y(_05408_));
 sky130_fd_sc_hd__o2bb2ai_2 _27943_ (.A1_N(_05399_),
    .A2_N(_05407_),
    .B1(_05288_),
    .B2(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__nor2_4 _27944_ (.A(_05288_),
    .B(_05408_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand3_4 _27945_ (.A(_05407_),
    .B(_05399_),
    .C(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__buf_2 _27946_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05412_));
 sky130_fd_sc_hd__buf_6 _27947_ (.A(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_8 _27948_ (.A(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__buf_6 _27949_ (.A(_05214_),
    .X(_05415_));
 sky130_fd_sc_hd__nand2_2 _27950_ (.A(_05414_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__buf_4 _27951_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05417_));
 sky130_fd_sc_hd__buf_4 _27952_ (.A(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__nand2_2 _27953_ (.A(_19918_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__nor2_4 _27954_ (.A(_05416_),
    .B(_05419_),
    .Y(_05420_));
 sky130_vsdinv _27955_ (.A(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__nand2_1 _27956_ (.A(_05416_),
    .B(_05419_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand2_2 _27957_ (.A(_05421_),
    .B(_05422_),
    .Y(_05423_));
 sky130_vsdinv _27958_ (.A(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__nand3_4 _27959_ (.A(_05409_),
    .B(_05411_),
    .C(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _27960_ (.A(_05407_),
    .B(_05399_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _27961_ (.A(_05426_),
    .B(_05410_),
    .Y(_05427_));
 sky130_fd_sc_hd__nand3b_2 _27962_ (.A_N(_05410_),
    .B(_05407_),
    .C(_05399_),
    .Y(_05428_));
 sky130_fd_sc_hd__nand3_4 _27963_ (.A(_05427_),
    .B(_05423_),
    .C(_05428_),
    .Y(_05429_));
 sky130_vsdinv _27964_ (.A(_05345_),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _27965_ (.A(_05343_),
    .B(_05344_),
    .Y(_05431_));
 sky130_fd_sc_hd__o2bb2ai_4 _27966_ (.A1_N(_05425_),
    .A2_N(_05429_),
    .B1(_05430_),
    .B2(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a21oi_2 _27967_ (.A1(_05341_),
    .A2(_05342_),
    .B1(_05430_),
    .Y(_05433_));
 sky130_fd_sc_hd__o2111ai_4 _27968_ (.A1(_05342_),
    .A2(_05341_),
    .B1(_05433_),
    .C1(_05425_),
    .D1(_05429_),
    .Y(_05434_));
 sky130_vsdinv _27969_ (.A(_05336_),
    .Y(_05435_));
 sky130_fd_sc_hd__and3_1 _27970_ (.A(_05327_),
    .B(_05255_),
    .C(_05280_),
    .X(_05436_));
 sky130_fd_sc_hd__or2_4 _27971_ (.A(_05435_),
    .B(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__a21o_1 _27972_ (.A1(_05432_),
    .A2(_05434_),
    .B1(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__nand3_4 _27973_ (.A(_05432_),
    .B(_05434_),
    .C(_05437_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand3_1 _27974_ (.A(_05363_),
    .B(_05438_),
    .C(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__nor3b_1 _27975_ (.A(_05362_),
    .B(_05360_),
    .C_N(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__nor2_2 _27976_ (.A(_05357_),
    .B(_05350_),
    .Y(_05442_));
 sky130_fd_sc_hd__a21oi_4 _27977_ (.A1(_05432_),
    .A2(_05434_),
    .B1(_05437_),
    .Y(_05443_));
 sky130_fd_sc_hd__o211a_4 _27978_ (.A1(_05435_),
    .A2(_05436_),
    .B1(_05434_),
    .C1(_05432_),
    .X(_05444_));
 sky130_fd_sc_hd__o22ai_2 _27979_ (.A1(_05351_),
    .A2(_05442_),
    .B1(_05443_),
    .B2(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o2bb2ai_1 _27980_ (.A1_N(_05440_),
    .A2_N(_05445_),
    .B1(_05362_),
    .B2(_05360_),
    .Y(_05446_));
 sky130_fd_sc_hd__a21boi_1 _27981_ (.A1(_05441_),
    .A2(_05445_),
    .B1_N(_05446_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21bo_1 _27982_ (.A1(_05397_),
    .A2(_05385_),
    .B1_N(_05381_),
    .X(_05447_));
 sky130_fd_sc_hd__nor2_4 _27983_ (.A(_05373_),
    .B(_05368_),
    .Y(_05448_));
 sky130_fd_sc_hd__nand2_4 _27984_ (.A(_05366_),
    .B(_05251_),
    .Y(_05449_));
 sky130_fd_sc_hd__buf_6 _27985_ (.A(_05227_),
    .X(_05450_));
 sky130_fd_sc_hd__buf_6 _27986_ (.A(_20167_),
    .X(_05451_));
 sky130_fd_sc_hd__nand3b_4 _27987_ (.A_N(_05449_),
    .B(_05450_),
    .C(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__buf_4 _27988_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05453_));
 sky130_fd_sc_hd__buf_6 _27989_ (.A(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__and2_2 _27990_ (.A(net469),
    .B(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__buf_4 _27991_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05456_));
 sky130_fd_sc_hd__nand2_4 _27992_ (.A(_05302_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__nand2_4 _27993_ (.A(_05449_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__nand3_4 _27994_ (.A(_05452_),
    .B(_05455_),
    .C(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__buf_6 _27995_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05460_));
 sky130_fd_sc_hd__a22oi_4 _27996_ (.A1(_05376_),
    .A2(_05176_),
    .B1(_05211_),
    .B2(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__nor2_4 _27997_ (.A(_05449_),
    .B(_05457_),
    .Y(_05462_));
 sky130_fd_sc_hd__buf_6 _27998_ (.A(_20151_),
    .X(_05463_));
 sky130_fd_sc_hd__nand2_4 _27999_ (.A(_19937_),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__o21ai_2 _28000_ (.A1(_05461_),
    .A2(_05462_),
    .B1(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__o211ai_4 _28001_ (.A1(_05371_),
    .A2(_05448_),
    .B1(_05459_),
    .C1(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21oi_2 _28002_ (.A1(_05378_),
    .A2(_05375_),
    .B1(_05371_),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_2 _28003_ (.A1(_05461_),
    .A2(_05462_),
    .B1(_05455_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand3_2 _28004_ (.A(_05452_),
    .B(_05464_),
    .C(_05458_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand3_4 _28005_ (.A(_05467_),
    .B(_05468_),
    .C(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_1 _28006_ (.A(_05466_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__buf_6 _28007_ (.A(_20154_),
    .X(_05472_));
 sky130_fd_sc_hd__nand2_2 _28008_ (.A(_05241_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__buf_6 _28009_ (.A(_05308_),
    .X(_05474_));
 sky130_fd_sc_hd__nand3_4 _28010_ (.A(_05473_),
    .B(_05282_),
    .C(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_2 _28011_ (.A(_05235_),
    .B(_05308_),
    .Y(_05476_));
 sky130_fd_sc_hd__buf_6 _28012_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05477_));
 sky130_fd_sc_hd__nand3_4 _28013_ (.A(_05476_),
    .B(_05477_),
    .C(_20156_),
    .Y(_05478_));
 sky130_fd_sc_hd__a21oi_1 _28014_ (.A1(_05475_),
    .A2(_05478_),
    .B1(_05154_),
    .Y(_05479_));
 sky130_fd_sc_hd__buf_4 _28015_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05480_));
 sky130_fd_sc_hd__buf_6 _28016_ (.A(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__nand2_1 _28017_ (.A(_05247_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__and3_1 _28018_ (.A(_05475_),
    .B(_05478_),
    .C(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__a21o_1 _28019_ (.A1(_05479_),
    .A2(_20163_),
    .B1(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__nand2_1 _28020_ (.A(_05471_),
    .B(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__a21oi_4 _28021_ (.A1(_05475_),
    .A2(_05478_),
    .B1(_05482_),
    .Y(_05486_));
 sky130_fd_sc_hd__nor2_4 _28022_ (.A(_05486_),
    .B(_05483_),
    .Y(_05487_));
 sky130_fd_sc_hd__nand3_2 _28023_ (.A(_05487_),
    .B(_05466_),
    .C(_05470_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand3_4 _28024_ (.A(_05447_),
    .B(_05485_),
    .C(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__a21boi_2 _28025_ (.A1(_05397_),
    .A2(_05385_),
    .B1_N(_05381_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_1 _28026_ (.A(_05471_),
    .B(_05487_),
    .Y(_05491_));
 sky130_fd_sc_hd__nand3_2 _28027_ (.A(_05484_),
    .B(_05470_),
    .C(_05466_),
    .Y(_05492_));
 sky130_fd_sc_hd__nand3_4 _28028_ (.A(_05490_),
    .B(_05491_),
    .C(_05492_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _28029_ (.A(_05489_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__o21ba_1 _28030_ (.A1(_05386_),
    .A2(_05390_),
    .B1_N(_05393_),
    .X(_05495_));
 sky130_fd_sc_hd__nand2_2 _28031_ (.A(_05494_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand3b_4 _28032_ (.A_N(_05495_),
    .B(_05489_),
    .C(_05493_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand2_1 _28033_ (.A(_05496_),
    .B(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__clkbuf_8 _28034_ (.A(_19914_),
    .X(_05499_));
 sky130_fd_sc_hd__nand2_4 _28035_ (.A(_05499_),
    .B(_05417_),
    .Y(_05500_));
 sky130_fd_sc_hd__buf_4 _28036_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05501_));
 sky130_fd_sc_hd__buf_4 _28037_ (.A(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__nand2_4 _28038_ (.A(net468),
    .B(_04838_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor2_4 _28039_ (.A(_05500_),
    .B(_05503_),
    .Y(_05504_));
 sky130_vsdinv _28040_ (.A(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__buf_6 _28041_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05506_));
 sky130_fd_sc_hd__nand2_2 _28042_ (.A(_05506_),
    .B(_05143_),
    .Y(_05507_));
 sky130_vsdinv _28043_ (.A(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__nand2_4 _28044_ (.A(_05500_),
    .B(_05503_),
    .Y(_05509_));
 sky130_fd_sc_hd__nand3_4 _28045_ (.A(_05505_),
    .B(_05508_),
    .C(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__buf_6 _28046_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05511_));
 sky130_fd_sc_hd__buf_1 _28047_ (.A(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__a22oi_4 _28048_ (.A1(net467),
    .A2(_05230_),
    .B1(_05414_),
    .B2(_05418_),
    .Y(_05513_));
 sky130_fd_sc_hd__o21ai_2 _28049_ (.A1(_05513_),
    .A2(_05504_),
    .B1(_05507_),
    .Y(_05514_));
 sky130_fd_sc_hd__a21o_1 _28050_ (.A1(_05510_),
    .A2(_05514_),
    .B1(_05420_),
    .X(_05515_));
 sky130_fd_sc_hd__nand3_4 _28051_ (.A(_05510_),
    .B(_05420_),
    .C(_05514_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_2 _28052_ (.A(_05515_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_4 _28053_ (.A(_05498_),
    .B(_05517_),
    .Y(_05518_));
 sky130_vsdinv _28054_ (.A(_05517_),
    .Y(_05519_));
 sky130_fd_sc_hd__nand3_2 _28055_ (.A(_05496_),
    .B(_05497_),
    .C(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__buf_6 _28056_ (.A(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__nand2_4 _28057_ (.A(_05518_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_4 _28058_ (.A(_05522_),
    .B(_05425_),
    .Y(_05523_));
 sky130_fd_sc_hd__and3_2 _28059_ (.A(_05409_),
    .B(_05411_),
    .C(_05424_),
    .X(_05524_));
 sky130_fd_sc_hd__nand3_4 _28060_ (.A(_05518_),
    .B(_05524_),
    .C(_05521_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_2 _28061_ (.A(_05523_),
    .B(_05525_),
    .Y(_05526_));
 sky130_vsdinv _28062_ (.A(_05399_),
    .Y(_05527_));
 sky130_fd_sc_hd__and2_1 _28063_ (.A(_05407_),
    .B(_05410_),
    .X(_05528_));
 sky130_fd_sc_hd__nor2_2 _28064_ (.A(_05346_),
    .B(_05524_),
    .Y(_05529_));
 sky130_fd_sc_hd__o211ai_4 _28065_ (.A1(_05527_),
    .A2(_05528_),
    .B1(_05429_),
    .C1(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_2 _28066_ (.A(_05527_),
    .B(_05528_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_4 _28067_ (.A(_05434_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand3_4 _28068_ (.A(_05526_),
    .B(_05530_),
    .C(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand2_2 _28069_ (.A(_05530_),
    .B(_05532_),
    .Y(_05534_));
 sky130_fd_sc_hd__nand3_4 _28070_ (.A(_05534_),
    .B(_05525_),
    .C(_05523_),
    .Y(_05535_));
 sky130_fd_sc_hd__o2111ai_4 _28071_ (.A1(_05351_),
    .A2(_05444_),
    .B1(_05438_),
    .C1(_05533_),
    .D1(_05535_),
    .Y(_05536_));
 sky130_vsdinv _28072_ (.A(_05520_),
    .Y(_05537_));
 sky130_fd_sc_hd__nand2_1 _28073_ (.A(_05518_),
    .B(_05524_),
    .Y(_05538_));
 sky130_fd_sc_hd__o2111ai_4 _28074_ (.A1(_05537_),
    .A2(_05538_),
    .B1(_05532_),
    .C1(_05523_),
    .D1(_05530_),
    .Y(_05539_));
 sky130_fd_sc_hd__nand2_1 _28075_ (.A(_05534_),
    .B(_05526_),
    .Y(_05540_));
 sky130_fd_sc_hd__o2111ai_4 _28076_ (.A1(_05355_),
    .A2(_05443_),
    .B1(_05439_),
    .C1(_05539_),
    .D1(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_2 _28077_ (.A(_05536_),
    .B(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__and3_1 _28078_ (.A(_05442_),
    .B(_05355_),
    .C(_05439_),
    .X(_05543_));
 sky130_fd_sc_hd__nand2_1 _28079_ (.A(_05543_),
    .B(_05438_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2_2 _28080_ (.A(_05446_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__xor2_1 _28081_ (.A(_05542_),
    .B(_05545_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_4 _28082_ (.A(_05535_),
    .B(_05533_),
    .Y(_05546_));
 sky130_fd_sc_hd__and3_1 _28083_ (.A(_05438_),
    .B(_05351_),
    .C(_05439_),
    .X(_05547_));
 sky130_fd_sc_hd__a22oi_4 _28084_ (.A1(_05546_),
    .A2(_05547_),
    .B1(_05545_),
    .B2(_05542_),
    .Y(_05548_));
 sky130_fd_sc_hd__buf_6 _28085_ (.A(_05243_),
    .X(_05549_));
 sky130_fd_sc_hd__a22oi_4 _28086_ (.A1(_05311_),
    .A2(_05549_),
    .B1(_05367_),
    .B2(_05388_),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_4 _28087_ (.A(_05227_),
    .B(_05251_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_4 _28088_ (.A(_19924_),
    .B(_05289_),
    .Y(_05552_));
 sky130_fd_sc_hd__nor2_4 _28089_ (.A(_05551_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__buf_4 _28090_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05554_));
 sky130_fd_sc_hd__buf_6 _28091_ (.A(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__nand2_4 _28092_ (.A(_05307_),
    .B(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__o21ai_4 _28093_ (.A1(_05550_),
    .A2(_05553_),
    .B1(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__buf_6 _28094_ (.A(_05366_),
    .X(_05558_));
 sky130_fd_sc_hd__nand3b_4 _28095_ (.A_N(_05551_),
    .B(_05558_),
    .C(_05286_),
    .Y(_05559_));
 sky130_vsdinv _28096_ (.A(_05556_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_4 _28097_ (.A(_05551_),
    .B(_05552_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand3_4 _28098_ (.A(_05559_),
    .B(_05560_),
    .C(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__o21ai_2 _28099_ (.A1(_05464_),
    .A2(_05461_),
    .B1(_05452_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand3_4 _28100_ (.A(_05557_),
    .B(_05562_),
    .C(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_2 _28101_ (.A1(_05550_),
    .A2(_05553_),
    .B1(_05560_),
    .Y(_05565_));
 sky130_fd_sc_hd__nand3_2 _28102_ (.A(_05559_),
    .B(_05556_),
    .C(_05561_),
    .Y(_05566_));
 sky130_fd_sc_hd__a21oi_2 _28103_ (.A1(_05458_),
    .A2(_05455_),
    .B1(_05462_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand3_4 _28104_ (.A(_05565_),
    .B(_05566_),
    .C(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand2_1 _28105_ (.A(_05564_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__buf_6 _28106_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05570_));
 sky130_fd_sc_hd__buf_4 _28107_ (.A(_05453_),
    .X(_05571_));
 sky130_fd_sc_hd__nand2_2 _28108_ (.A(_05570_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__buf_4 _28109_ (.A(_20155_),
    .X(_05573_));
 sky130_fd_sc_hd__nand3_4 _28110_ (.A(_05572_),
    .B(_19931_),
    .C(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand2_2 _28111_ (.A(_05387_),
    .B(_05472_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand3_4 _28112_ (.A(_05575_),
    .B(_05242_),
    .C(_20152_),
    .Y(_05576_));
 sky130_fd_sc_hd__buf_4 _28113_ (.A(_20158_),
    .X(_05577_));
 sky130_fd_sc_hd__nand2_1 _28114_ (.A(_05247_),
    .B(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__a21oi_4 _28115_ (.A1(_05574_),
    .A2(_05576_),
    .B1(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__buf_6 _28116_ (.A(_05295_),
    .X(_05580_));
 sky130_fd_sc_hd__o211a_2 _28117_ (.A1(_05186_),
    .A2(_05580_),
    .B1(_05574_),
    .C1(_05576_),
    .X(_05581_));
 sky130_fd_sc_hd__nor2_4 _28118_ (.A(_05579_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__nand2_1 _28119_ (.A(_05569_),
    .B(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21a_1 _28120_ (.A1(_05461_),
    .A2(_05462_),
    .B1(_05464_),
    .X(_05584_));
 sky130_fd_sc_hd__o21ai_2 _28121_ (.A1(_05371_),
    .A2(_05448_),
    .B1(_05459_),
    .Y(_05585_));
 sky130_fd_sc_hd__a2bb2oi_2 _28122_ (.A1_N(_05584_),
    .A2_N(_05585_),
    .B1(_05470_),
    .B2(_05487_),
    .Y(_05586_));
 sky130_fd_sc_hd__o211ai_4 _28123_ (.A1(_05579_),
    .A2(_05581_),
    .B1(_05564_),
    .C1(_05568_),
    .Y(_05587_));
 sky130_fd_sc_hd__nand3_4 _28124_ (.A(_05583_),
    .B(_05586_),
    .C(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__o2bb2ai_2 _28125_ (.A1_N(_05470_),
    .A2_N(_05487_),
    .B1(_05584_),
    .B2(_05585_),
    .Y(_05589_));
 sky130_fd_sc_hd__o2bb2ai_1 _28126_ (.A1_N(_05564_),
    .A2_N(_05568_),
    .B1(_05579_),
    .B2(_05581_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand3_2 _28127_ (.A(_05582_),
    .B(_05564_),
    .C(_05568_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand3_4 _28128_ (.A(_05589_),
    .B(_05590_),
    .C(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__nor2_4 _28129_ (.A(_05476_),
    .B(_05473_),
    .Y(_05593_));
 sky130_fd_sc_hd__or2_2 _28130_ (.A(_05593_),
    .B(_05486_),
    .X(_05594_));
 sky130_fd_sc_hd__a21o_1 _28131_ (.A1(_05588_),
    .A2(_05592_),
    .B1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__nand3_2 _28132_ (.A(_05588_),
    .B(_05592_),
    .C(_05594_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand2_4 _28133_ (.A(_05511_),
    .B(_20173_),
    .Y(_05597_));
 sky130_fd_sc_hd__buf_6 _28134_ (.A(_05412_),
    .X(_05598_));
 sky130_fd_sc_hd__nand2_4 _28135_ (.A(_05598_),
    .B(_05178_),
    .Y(_05599_));
 sky130_fd_sc_hd__or2_2 _28136_ (.A(_05597_),
    .B(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__buf_6 _28137_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05601_));
 sky130_fd_sc_hd__buf_6 _28138_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05602_));
 sky130_fd_sc_hd__nand2_2 _28139_ (.A(_05601_),
    .B(_05602_),
    .Y(_05603_));
 sky130_vsdinv _28140_ (.A(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__nand2_4 _28141_ (.A(_05597_),
    .B(_05599_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand3_4 _28142_ (.A(_05600_),
    .B(_05604_),
    .C(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__a21o_1 _28143_ (.A1(_05508_),
    .A2(_05509_),
    .B1(_05504_),
    .X(_05607_));
 sky130_fd_sc_hd__buf_8 _28144_ (.A(_05598_),
    .X(_05608_));
 sky130_fd_sc_hd__a22oi_4 _28145_ (.A1(_19912_),
    .A2(_20174_),
    .B1(_05608_),
    .B2(_05179_),
    .Y(_05609_));
 sky130_fd_sc_hd__nor2_4 _28146_ (.A(_05597_),
    .B(_05599_),
    .Y(_05610_));
 sky130_fd_sc_hd__o21ai_2 _28147_ (.A1(_05609_),
    .A2(_05610_),
    .B1(_05603_),
    .Y(_05611_));
 sky130_fd_sc_hd__nand3_4 _28148_ (.A(_05606_),
    .B(_05607_),
    .C(_05611_),
    .Y(_05612_));
 sky130_vsdinv _28149_ (.A(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand2_1 _28150_ (.A(_05514_),
    .B(_05420_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand3_4 _28151_ (.A(_05600_),
    .B(_05603_),
    .C(_05605_),
    .Y(_05615_));
 sky130_fd_sc_hd__a21oi_4 _28152_ (.A1(_05508_),
    .A2(_05509_),
    .B1(_05504_),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_2 _28153_ (.A1(_05609_),
    .A2(_05610_),
    .B1(_05604_),
    .Y(_05617_));
 sky130_fd_sc_hd__nand3_4 _28154_ (.A(_05615_),
    .B(_05616_),
    .C(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand3b_4 _28155_ (.A_N(_05614_),
    .B(_05618_),
    .C(_05510_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand2_1 _28156_ (.A(_05612_),
    .B(_05618_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _28157_ (.A(_05620_),
    .B(_05516_),
    .Y(_05621_));
 sky130_fd_sc_hd__o21a_4 _28158_ (.A1(_05613_),
    .A2(_05619_),
    .B1(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__nand3_4 _28159_ (.A(_05595_),
    .B(_05596_),
    .C(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__o2bb2ai_2 _28160_ (.A1_N(_05592_),
    .A2_N(_05588_),
    .B1(_05593_),
    .B2(_05486_),
    .Y(_05624_));
 sky130_fd_sc_hd__or2_2 _28161_ (.A(_05516_),
    .B(_05620_),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _28162_ (.A(_05625_),
    .B(_05621_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand3b_4 _28163_ (.A_N(_05594_),
    .B(_05588_),
    .C(_05592_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand3_4 _28164_ (.A(_05624_),
    .B(_05626_),
    .C(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__a32oi_4 _28165_ (.A1(_05496_),
    .A2(_05497_),
    .A3(_05519_),
    .B1(_05623_),
    .B2(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__nand2_4 _28166_ (.A(_05623_),
    .B(_05628_),
    .Y(_05630_));
 sky130_fd_sc_hd__nor2_8 _28167_ (.A(_05521_),
    .B(_05630_),
    .Y(_05631_));
 sky130_vsdinv _28168_ (.A(_19908_),
    .Y(_05632_));
 sky130_fd_sc_hd__buf_4 _28169_ (.A(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__nor2_2 _28170_ (.A(net448),
    .B(_04841_),
    .Y(_05634_));
 sky130_vsdinv _28171_ (.A(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ai_4 _28172_ (.A1(_05629_),
    .A2(_05631_),
    .B1(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__a21oi_4 _28173_ (.A1(_05630_),
    .A2(_05521_),
    .B1(_05635_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand3_4 _28174_ (.A(_05537_),
    .B(_05623_),
    .C(_05628_),
    .Y(_05638_));
 sky130_fd_sc_hd__nand2_4 _28175_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a21o_1 _28176_ (.A1(_05489_),
    .A2(_05497_),
    .B1(_05525_),
    .X(_05640_));
 sky130_fd_sc_hd__nand2_1 _28177_ (.A(_05497_),
    .B(_05489_),
    .Y(_05641_));
 sky130_fd_sc_hd__a31o_2 _28178_ (.A1(_05518_),
    .A2(_05524_),
    .A3(_05521_),
    .B1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__a22oi_2 _28179_ (.A1(_05636_),
    .A2(_05639_),
    .B1(_05640_),
    .B2(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__and4_1 _28180_ (.A(_05640_),
    .B(_05636_),
    .C(_05639_),
    .D(_05642_),
    .X(_05644_));
 sky130_fd_sc_hd__nor2_1 _28181_ (.A(_05531_),
    .B(_05434_),
    .Y(_05645_));
 sky130_fd_sc_hd__a31o_1 _28182_ (.A1(_05523_),
    .A2(_05525_),
    .A3(_05532_),
    .B1(_05645_),
    .X(_05646_));
 sky130_vsdinv _28183_ (.A(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_2 _28184_ (.A1(_05643_),
    .A2(_05644_),
    .B1(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__a22o_1 _28185_ (.A1(_05636_),
    .A2(_05639_),
    .B1(_05640_),
    .B2(_05642_),
    .X(_05649_));
 sky130_fd_sc_hd__nand2_2 _28186_ (.A(_05524_),
    .B(_05641_),
    .Y(_05650_));
 sky130_fd_sc_hd__o2111ai_4 _28187_ (.A1(_05522_),
    .A2(_05650_),
    .B1(_05642_),
    .C1(_05639_),
    .D1(_05636_),
    .Y(_05651_));
 sky130_fd_sc_hd__nand3_4 _28188_ (.A(_05649_),
    .B(_05646_),
    .C(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__a22oi_4 _28189_ (.A1(_05444_),
    .A2(_05546_),
    .B1(_05648_),
    .B2(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__a31o_1 _28190_ (.A1(_05444_),
    .A2(_05546_),
    .A3(_05648_),
    .B1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__xor2_1 _28191_ (.A(_05548_),
    .B(_05654_),
    .X(_02686_));
 sky130_vsdinv _28192_ (.A(_05652_),
    .Y(_05655_));
 sky130_fd_sc_hd__buf_4 _28193_ (.A(\pcpi_mul.rs2[10] ),
    .X(_05656_));
 sky130_fd_sc_hd__buf_8 _28194_ (.A(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__nand2_4 _28195_ (.A(_05657_),
    .B(_20177_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_4 _28196_ (.A(_19909_),
    .B(_05146_),
    .Y(_05659_));
 sky130_fd_sc_hd__nor2_8 _28197_ (.A(_05658_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand2_1 _28198_ (.A(_05658_),
    .B(_05659_),
    .Y(_05661_));
 sky130_vsdinv _28199_ (.A(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__nand2_2 _28200_ (.A(_05624_),
    .B(_05627_),
    .Y(_05663_));
 sky130_fd_sc_hd__buf_6 _28201_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05664_));
 sky130_fd_sc_hd__buf_6 _28202_ (.A(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__a22oi_4 _28203_ (.A1(_05450_),
    .A2(_20162_),
    .B1(_05558_),
    .B2(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_2 _28204_ (.A(_05302_),
    .B(_05480_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_2 _28205_ (.A(_05211_),
    .B(_20158_),
    .Y(_05668_));
 sky130_fd_sc_hd__nor2_2 _28206_ (.A(_05667_),
    .B(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__buf_4 _28207_ (.A(_20144_),
    .X(_05670_));
 sky130_fd_sc_hd__nand2_2 _28208_ (.A(_05307_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__clkbuf_2 _28209_ (.A(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__o21bai_2 _28210_ (.A1(_05666_),
    .A2(_05669_),
    .B1_N(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__buf_6 _28211_ (.A(_05211_),
    .X(_05674_));
 sky130_fd_sc_hd__buf_4 _28212_ (.A(_05391_),
    .X(_05675_));
 sky130_fd_sc_hd__nand3b_4 _28213_ (.A_N(_05667_),
    .B(_05674_),
    .C(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_2 _28214_ (.A(_05667_),
    .B(_05668_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand3_2 _28215_ (.A(_05676_),
    .B(_05677_),
    .C(_05672_),
    .Y(_05678_));
 sky130_fd_sc_hd__o21ai_1 _28216_ (.A1(_05551_),
    .A2(_05552_),
    .B1(_05556_),
    .Y(_05679_));
 sky130_fd_sc_hd__nand2_1 _28217_ (.A(_05679_),
    .B(_05561_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand3_4 _28218_ (.A(_05673_),
    .B(_05678_),
    .C(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__o21ai_2 _28219_ (.A1(_05666_),
    .A2(_05669_),
    .B1(_05672_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21ai_4 _28220_ (.A1(_05556_),
    .A2(_05550_),
    .B1(_05559_),
    .Y(_05683_));
 sky130_fd_sc_hd__buf_6 _28221_ (.A(_05308_),
    .X(_05684_));
 sky130_fd_sc_hd__a41oi_2 _28222_ (.A1(_19920_),
    .A2(_05298_),
    .A3(_05684_),
    .A4(_05286_),
    .B1(_05671_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand2_2 _28223_ (.A(_05685_),
    .B(_05677_),
    .Y(_05686_));
 sky130_fd_sc_hd__nand3_4 _28224_ (.A(_05682_),
    .B(_05683_),
    .C(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__a22oi_4 _28225_ (.A1(_05282_),
    .A2(_05463_),
    .B1(_05284_),
    .B2(_20149_),
    .Y(_05688_));
 sky130_fd_sc_hd__buf_6 _28226_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05689_));
 sky130_fd_sc_hd__nand2_8 _28227_ (.A(_05689_),
    .B(_20151_),
    .Y(_05690_));
 sky130_fd_sc_hd__nor2_8 _28228_ (.A(_05129_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__buf_6 _28229_ (.A(_19927_),
    .X(_05692_));
 sky130_fd_sc_hd__buf_4 _28230_ (.A(_05472_),
    .X(_05693_));
 sky130_fd_sc_hd__nand2_2 _28231_ (.A(_05692_),
    .B(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_2 _28232_ (.A1(_05688_),
    .A2(_05691_),
    .B1(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__buf_6 _28233_ (.A(_20154_),
    .X(_05696_));
 sky130_fd_sc_hd__buf_6 _28234_ (.A(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__buf_4 _28235_ (.A(_05453_),
    .X(_05698_));
 sky130_fd_sc_hd__buf_6 _28236_ (.A(_05554_),
    .X(_05699_));
 sky130_fd_sc_hd__a22o_1 _28237_ (.A1(_05173_),
    .A2(_05698_),
    .B1(_05477_),
    .B2(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__o2111ai_4 _28238_ (.A1(_05130_),
    .A2(_05690_),
    .B1(_05692_),
    .C1(_05697_),
    .D1(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand2_4 _28239_ (.A(_05695_),
    .B(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__a21o_1 _28240_ (.A1(_05681_),
    .A2(_05687_),
    .B1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_1 _28241_ (.A(_05458_),
    .B(_05455_),
    .Y(_05704_));
 sky130_fd_sc_hd__a32oi_4 _28242_ (.A1(_05559_),
    .A2(_05560_),
    .A3(_05561_),
    .B1(_05452_),
    .B2(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__a22oi_4 _28243_ (.A1(_05705_),
    .A2(_05557_),
    .B1(_05582_),
    .B2(_05568_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand3_2 _28244_ (.A(_05681_),
    .B(_05687_),
    .C(_05702_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand3_4 _28245_ (.A(_05703_),
    .B(_05706_),
    .C(_05707_),
    .Y(_05708_));
 sky130_vsdinv _28246_ (.A(_05557_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand2_1 _28247_ (.A(_05562_),
    .B(_05563_),
    .Y(_05710_));
 sky130_fd_sc_hd__o2bb2ai_2 _28248_ (.A1_N(_05568_),
    .A2_N(_05582_),
    .B1(_05709_),
    .B2(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__nor3_4 _28249_ (.A(_05694_),
    .B(_05688_),
    .C(_05691_),
    .Y(_05712_));
 sky130_fd_sc_hd__o21a_1 _28250_ (.A1(_05688_),
    .A2(_05691_),
    .B1(_05694_),
    .X(_05713_));
 sky130_fd_sc_hd__o2bb2ai_2 _28251_ (.A1_N(_05681_),
    .A2_N(_05687_),
    .B1(_05712_),
    .B2(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__nand3b_4 _28252_ (.A_N(_05702_),
    .B(_05681_),
    .C(_05687_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand3_4 _28253_ (.A(_05711_),
    .B(_05714_),
    .C(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__nand2_1 _28254_ (.A(_05708_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__nor2_4 _28255_ (.A(_05575_),
    .B(_05572_),
    .Y(_05718_));
 sky130_fd_sc_hd__nor2_2 _28256_ (.A(_05718_),
    .B(_05579_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand2_2 _28257_ (.A(_05717_),
    .B(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__nand2_1 _28258_ (.A(_05606_),
    .B(_05611_),
    .Y(_05721_));
 sky130_fd_sc_hd__buf_6 _28259_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05722_));
 sky130_fd_sc_hd__nand2_4 _28260_ (.A(_05722_),
    .B(_20170_),
    .Y(_05723_));
 sky130_fd_sc_hd__buf_6 _28261_ (.A(_05412_),
    .X(_05724_));
 sky130_fd_sc_hd__nand2_4 _28262_ (.A(_05724_),
    .B(_05456_),
    .Y(_05725_));
 sky130_fd_sc_hd__nor2_8 _28263_ (.A(_05723_),
    .B(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__and2_2 _28264_ (.A(_05723_),
    .B(_05725_),
    .X(_05727_));
 sky130_fd_sc_hd__nand2_2 _28265_ (.A(_05601_),
    .B(_05237_),
    .Y(_05728_));
 sky130_vsdinv _28266_ (.A(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__o21ai_2 _28267_ (.A1(_05726_),
    .A2(_05727_),
    .B1(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__or2_2 _28268_ (.A(_05723_),
    .B(_05725_),
    .X(_05731_));
 sky130_fd_sc_hd__nand2_2 _28269_ (.A(_05723_),
    .B(_05725_),
    .Y(_05732_));
 sky130_fd_sc_hd__nand3_2 _28270_ (.A(_05731_),
    .B(_05728_),
    .C(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__a21oi_2 _28271_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05610_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand3_4 _28272_ (.A(_05730_),
    .B(_05733_),
    .C(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__o21ai_4 _28273_ (.A1(_05726_),
    .A2(_05727_),
    .B1(_05728_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand3_4 _28274_ (.A(_05731_),
    .B(_05729_),
    .C(_05732_),
    .Y(_05737_));
 sky130_fd_sc_hd__a21o_2 _28275_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05610_),
    .X(_05738_));
 sky130_fd_sc_hd__nand3_4 _28276_ (.A(_05736_),
    .B(_05737_),
    .C(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__o2111ai_4 _28277_ (.A1(_05616_),
    .A2(_05721_),
    .B1(_05735_),
    .C1(_05739_),
    .D1(_05619_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_4 _28278_ (.A(_05739_),
    .B(_05735_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _28279_ (.A(_05516_),
    .B(_05612_),
    .Y(_05742_));
 sky130_fd_sc_hd__nand3_4 _28280_ (.A(_05741_),
    .B(_05742_),
    .C(_05618_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_4 _28281_ (.A(_05740_),
    .B(_05743_),
    .Y(_05744_));
 sky130_vsdinv _28282_ (.A(_05719_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand3_4 _28283_ (.A(_05708_),
    .B(_05716_),
    .C(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__nand3_2 _28284_ (.A(_05720_),
    .B(_05744_),
    .C(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__o2bb2ai_2 _28285_ (.A1_N(_05708_),
    .A2_N(_05716_),
    .B1(_05718_),
    .B2(_05579_),
    .Y(_05748_));
 sky130_fd_sc_hd__and2_1 _28286_ (.A(_05740_),
    .B(_05743_),
    .X(_05749_));
 sky130_fd_sc_hd__nand3_2 _28287_ (.A(_05708_),
    .B(_05716_),
    .C(_05719_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand3_4 _28288_ (.A(_05748_),
    .B(_05749_),
    .C(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__a22oi_4 _28289_ (.A1(_05663_),
    .A2(_05622_),
    .B1(_05747_),
    .B2(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__a21oi_4 _28290_ (.A1(_05708_),
    .A2(_05716_),
    .B1(_05745_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_4 _28291_ (.A(_05746_),
    .B(_05744_),
    .Y(_05754_));
 sky130_fd_sc_hd__o2111a_1 _28292_ (.A1(_05753_),
    .A2(_05754_),
    .B1(_05622_),
    .C1(_05663_),
    .D1(_05751_),
    .X(_05755_));
 sky130_fd_sc_hd__o22ai_4 _28293_ (.A1(_05660_),
    .A2(_05662_),
    .B1(_05752_),
    .B2(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21ai_2 _28294_ (.A1(_05753_),
    .A2(_05754_),
    .B1(_05751_),
    .Y(_05757_));
 sky130_fd_sc_hd__nand2_4 _28295_ (.A(_05757_),
    .B(_05623_),
    .Y(_05758_));
 sky130_fd_sc_hd__o2111ai_4 _28296_ (.A1(_05753_),
    .A2(_05754_),
    .B1(_05622_),
    .C1(_05663_),
    .D1(_05751_),
    .Y(_05759_));
 sky130_fd_sc_hd__buf_4 _28297_ (.A(_05759_),
    .X(_05760_));
 sky130_vsdinv _28298_ (.A(_05660_),
    .Y(_05761_));
 sky130_fd_sc_hd__nand2_2 _28299_ (.A(_05761_),
    .B(_05661_),
    .Y(_05762_));
 sky130_vsdinv _28300_ (.A(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand3_4 _28301_ (.A(_05758_),
    .B(_05760_),
    .C(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__a22oi_4 _28302_ (.A1(_05638_),
    .A2(_05637_),
    .B1(_05756_),
    .B2(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__a21oi_4 _28303_ (.A1(_05758_),
    .A2(_05760_),
    .B1(_05763_),
    .Y(_05766_));
 sky130_fd_sc_hd__nand3_2 _28304_ (.A(_05764_),
    .B(_05638_),
    .C(_05637_),
    .Y(_05767_));
 sky130_fd_sc_hd__nor2_4 _28305_ (.A(_05766_),
    .B(_05767_),
    .Y(_05768_));
 sky130_vsdinv _28306_ (.A(_05592_),
    .Y(_05769_));
 sky130_fd_sc_hd__and2_2 _28307_ (.A(_05588_),
    .B(_05594_),
    .X(_05770_));
 sky130_fd_sc_hd__nor2_8 _28308_ (.A(_05769_),
    .B(_05770_),
    .Y(_05771_));
 sky130_vsdinv _28309_ (.A(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__nor2_4 _28310_ (.A(_05772_),
    .B(_05631_),
    .Y(_05773_));
 sky130_fd_sc_hd__nor2_4 _28311_ (.A(_05771_),
    .B(_05638_),
    .Y(_05774_));
 sky130_fd_sc_hd__nor2_2 _28312_ (.A(_05773_),
    .B(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__o21ai_2 _28313_ (.A1(_05765_),
    .A2(_05768_),
    .B1(_05775_),
    .Y(_05776_));
 sky130_fd_sc_hd__nor2_2 _28314_ (.A(_05650_),
    .B(_05522_),
    .Y(_05777_));
 sky130_fd_sc_hd__a31oi_4 _28315_ (.A1(_05636_),
    .A2(_05639_),
    .A3(_05642_),
    .B1(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__and3_2 _28316_ (.A(_05758_),
    .B(_05759_),
    .C(_05763_),
    .X(_05779_));
 sky130_fd_sc_hd__o21ai_2 _28317_ (.A1(_05766_),
    .A2(_05779_),
    .B1(_05639_),
    .Y(_05780_));
 sky130_fd_sc_hd__o2111ai_4 _28318_ (.A1(_05521_),
    .A2(_05630_),
    .B1(_05637_),
    .C1(_05764_),
    .D1(_05756_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_1 _28319_ (.A(_05638_),
    .B(_05771_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand2_1 _28320_ (.A(_05631_),
    .B(_05772_),
    .Y(_05783_));
 sky130_fd_sc_hd__nand2_2 _28321_ (.A(_05782_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__nand3_2 _28322_ (.A(_05780_),
    .B(_05781_),
    .C(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand3_4 _28323_ (.A(_05776_),
    .B(_05778_),
    .C(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2_1 _28324_ (.A(_05649_),
    .B(_05651_),
    .Y(_05787_));
 sky130_fd_sc_hd__o22ai_4 _28325_ (.A1(_05773_),
    .A2(_05774_),
    .B1(_05765_),
    .B2(_05768_),
    .Y(_05788_));
 sky130_fd_sc_hd__nand3_2 _28326_ (.A(_05780_),
    .B(_05775_),
    .C(_05781_),
    .Y(_05789_));
 sky130_fd_sc_hd__nand2_1 _28327_ (.A(_05651_),
    .B(_05640_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand3_4 _28328_ (.A(_05788_),
    .B(_05789_),
    .C(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__a2bb2oi_2 _28329_ (.A1_N(_05787_),
    .A2_N(_05647_),
    .B1(_05791_),
    .B2(_05786_),
    .Y(_05792_));
 sky130_fd_sc_hd__a21oi_4 _28330_ (.A1(_05655_),
    .A2(_05786_),
    .B1(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_1 _28331_ (.A(_05546_),
    .B(_05444_),
    .Y(_05794_));
 sky130_vsdinv _28332_ (.A(_05648_),
    .Y(_05795_));
 sky130_fd_sc_hd__o22ai_4 _28333_ (.A1(_05794_),
    .A2(_05795_),
    .B1(_05653_),
    .B2(_05548_),
    .Y(_05796_));
 sky130_fd_sc_hd__xor2_1 _28334_ (.A(_05793_),
    .B(_05796_),
    .X(_02629_));
 sky130_fd_sc_hd__buf_6 _28335_ (.A(_05302_),
    .X(_05797_));
 sky130_fd_sc_hd__a22oi_4 _28336_ (.A1(_05797_),
    .A2(_05684_),
    .B1(_19925_),
    .B2(_05573_),
    .Y(_05798_));
 sky130_fd_sc_hd__buf_6 _28337_ (.A(_20154_),
    .X(_05799_));
 sky130_fd_sc_hd__and4_4 _28338_ (.A(_05450_),
    .B(_05312_),
    .C(_05799_),
    .D(_05389_),
    .X(_05800_));
 sky130_fd_sc_hd__nand2_2 _28339_ (.A(_19937_),
    .B(_20142_),
    .Y(_05801_));
 sky130_vsdinv _28340_ (.A(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21ai_2 _28341_ (.A1(_05798_),
    .A2(_05800_),
    .B1(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand2_1 _28342_ (.A(_05797_),
    .B(_05474_),
    .Y(_05804_));
 sky130_fd_sc_hd__buf_6 _28343_ (.A(_05558_),
    .X(_05805_));
 sky130_fd_sc_hd__nand3b_4 _28344_ (.A_N(_05804_),
    .B(_05805_),
    .C(_20157_),
    .Y(_05806_));
 sky130_fd_sc_hd__a22o_2 _28345_ (.A1(_05797_),
    .A2(_05684_),
    .B1(_05298_),
    .B2(_05573_),
    .X(_05807_));
 sky130_fd_sc_hd__nand3_2 _28346_ (.A(_05806_),
    .B(_05807_),
    .C(_05801_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ai_1 _28347_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05672_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _28348_ (.A(_05809_),
    .B(_05677_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand3_4 _28349_ (.A(_05803_),
    .B(_05808_),
    .C(_05810_),
    .Y(_05811_));
 sky130_vsdinv _28350_ (.A(_20141_),
    .Y(_05812_));
 sky130_fd_sc_hd__clkbuf_8 _28351_ (.A(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__o22ai_4 _28352_ (.A1(net470),
    .A2(_05813_),
    .B1(_05798_),
    .B2(_05800_),
    .Y(_05814_));
 sky130_fd_sc_hd__o21ai_2 _28353_ (.A1(_05672_),
    .A2(_05666_),
    .B1(_05676_),
    .Y(_05815_));
 sky130_fd_sc_hd__buf_6 _28354_ (.A(_05376_),
    .X(_05816_));
 sky130_fd_sc_hd__a41oi_1 _28355_ (.A1(_05816_),
    .A2(_05674_),
    .A3(_05693_),
    .A4(_05675_),
    .B1(_05801_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _28356_ (.A(_05817_),
    .B(_05807_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand3_4 _28357_ (.A(_05814_),
    .B(_05815_),
    .C(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__buf_8 _28358_ (.A(_05555_),
    .X(_05820_));
 sky130_fd_sc_hd__buf_4 _28359_ (.A(_05241_),
    .X(_05821_));
 sky130_fd_sc_hd__buf_6 _28360_ (.A(_20144_),
    .X(_05822_));
 sky130_fd_sc_hd__buf_8 _28361_ (.A(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__a22oi_4 _28362_ (.A1(_05236_),
    .A2(_05820_),
    .B1(_05821_),
    .B2(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__clkbuf_4 _28363_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_8 _28364_ (.A(_05825_),
    .X(_05826_));
 sky130_fd_sc_hd__buf_8 _28365_ (.A(_05554_),
    .X(_05827_));
 sky130_fd_sc_hd__nand2_8 _28366_ (.A(_05826_),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__nor2_8 _28367_ (.A(_05130_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__buf_4 _28368_ (.A(_19927_),
    .X(_05830_));
 sky130_fd_sc_hd__buf_6 _28369_ (.A(_20151_),
    .X(_05831_));
 sky130_fd_sc_hd__buf_6 _28370_ (.A(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__nand2_1 _28371_ (.A(_05830_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__o21ai_1 _28372_ (.A1(_05824_),
    .A2(_05829_),
    .B1(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__buf_4 _28373_ (.A(_05670_),
    .X(_05835_));
 sky130_fd_sc_hd__a22o_1 _28374_ (.A1(_19931_),
    .A2(_20149_),
    .B1(_05242_),
    .B2(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__o2111ai_4 _28375_ (.A1(_05130_),
    .A2(_05828_),
    .B1(_19928_),
    .C1(_05832_),
    .D1(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_2 _28376_ (.A(_05834_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__a21o_1 _28377_ (.A1(_05811_),
    .A2(_05819_),
    .B1(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_1 _28378_ (.A(_05687_),
    .B(_05702_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _28379_ (.A(_05840_),
    .B(_05681_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand3_2 _28380_ (.A(_05811_),
    .B(_05819_),
    .C(_05838_),
    .Y(_05842_));
 sky130_fd_sc_hd__nand3_4 _28381_ (.A(_05839_),
    .B(_05841_),
    .C(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__o21a_1 _28382_ (.A1(_05666_),
    .A2(_05669_),
    .B1(_05672_),
    .X(_05844_));
 sky130_fd_sc_hd__nand2_1 _28383_ (.A(_05683_),
    .B(_05686_),
    .Y(_05845_));
 sky130_fd_sc_hd__a21oi_2 _28384_ (.A1(_05682_),
    .A2(_05686_),
    .B1(_05683_),
    .Y(_05846_));
 sky130_fd_sc_hd__o22ai_4 _28385_ (.A1(_05844_),
    .A2(_05845_),
    .B1(_05702_),
    .B2(_05846_),
    .Y(_05847_));
 sky130_vsdinv _28386_ (.A(_05837_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21a_1 _28387_ (.A1(_05824_),
    .A2(_05829_),
    .B1(_05833_),
    .X(_05849_));
 sky130_fd_sc_hd__o2bb2ai_2 _28388_ (.A1_N(_05819_),
    .A2_N(_05811_),
    .B1(_05848_),
    .B2(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__nand3b_2 _28389_ (.A_N(_05838_),
    .B(_05811_),
    .C(_05819_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand3_4 _28390_ (.A(_05847_),
    .B(_05850_),
    .C(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__nand2_1 _28391_ (.A(_05843_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__nor2_2 _28392_ (.A(_05691_),
    .B(_05712_),
    .Y(_05854_));
 sky130_fd_sc_hd__nand2_1 _28393_ (.A(_05853_),
    .B(_05854_),
    .Y(_05855_));
 sky130_vsdinv _28394_ (.A(_05854_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand3_2 _28395_ (.A(_05843_),
    .B(_05852_),
    .C(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__buf_6 _28396_ (.A(_19911_),
    .X(_05858_));
 sky130_fd_sc_hd__a22oi_4 _28397_ (.A1(_05858_),
    .A2(_05183_),
    .B1(_05414_),
    .B2(_05238_),
    .Y(_05859_));
 sky130_fd_sc_hd__nand2_8 _28398_ (.A(_05501_),
    .B(_19914_),
    .Y(_05860_));
 sky130_fd_sc_hd__buf_8 _28399_ (.A(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__nand2_1 _28400_ (.A(_05237_),
    .B(_05602_),
    .Y(_05862_));
 sky130_fd_sc_hd__buf_4 _28401_ (.A(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__nor2_2 _28402_ (.A(_05861_),
    .B(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__buf_6 _28403_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05865_));
 sky130_fd_sc_hd__buf_6 _28404_ (.A(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__clkbuf_8 _28405_ (.A(_05480_),
    .X(_05867_));
 sky130_fd_sc_hd__nand2_2 _28406_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_2 _28407_ (.A1(_05859_),
    .A2(_05864_),
    .B1(_05868_),
    .Y(_05869_));
 sky130_vsdinv _28408_ (.A(_05868_),
    .Y(_05870_));
 sky130_fd_sc_hd__a22o_2 _28409_ (.A1(net467),
    .A2(_05177_),
    .B1(_05608_),
    .B2(_05238_),
    .X(_05871_));
 sky130_fd_sc_hd__o211ai_4 _28410_ (.A1(_05861_),
    .A2(_05863_),
    .B1(_05870_),
    .C1(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand3_4 _28411_ (.A(_05869_),
    .B(_05660_),
    .C(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__o21ai_2 _28412_ (.A1(_05859_),
    .A2(_05864_),
    .B1(_05870_),
    .Y(_05874_));
 sky130_fd_sc_hd__o211ai_4 _28413_ (.A1(_05861_),
    .A2(_05863_),
    .B1(_05868_),
    .C1(_05871_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand3_4 _28414_ (.A(_05874_),
    .B(_05761_),
    .C(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__nor2_4 _28415_ (.A(_05729_),
    .B(_05726_),
    .Y(_05877_));
 sky130_fd_sc_hd__o2bb2ai_4 _28416_ (.A1_N(_05873_),
    .A2_N(_05876_),
    .B1(_05727_),
    .B2(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__nor2_2 _28417_ (.A(_05727_),
    .B(_05877_),
    .Y(_05879_));
 sky130_fd_sc_hd__nand3_4 _28418_ (.A(_05873_),
    .B(_05876_),
    .C(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__nand2_4 _28419_ (.A(_05878_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__a21oi_4 _28420_ (.A1(_05736_),
    .A2(_05737_),
    .B1(_05738_),
    .Y(_05882_));
 sky130_fd_sc_hd__o21ai_1 _28421_ (.A1(_05612_),
    .A2(_05882_),
    .B1(_05739_),
    .Y(_05883_));
 sky130_fd_sc_hd__nand2_1 _28422_ (.A(_05881_),
    .B(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__o2111ai_4 _28423_ (.A1(_05612_),
    .A2(_05882_),
    .B1(_05739_),
    .C1(_05880_),
    .D1(_05878_),
    .Y(_05885_));
 sky130_fd_sc_hd__nand2_1 _28424_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__nand3_4 _28425_ (.A(_05855_),
    .B(_05857_),
    .C(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__o2bb2ai_2 _28426_ (.A1_N(_05843_),
    .A2_N(_05852_),
    .B1(_05691_),
    .B2(_05712_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand3_2 _28427_ (.A(_05843_),
    .B(_05852_),
    .C(_05854_),
    .Y(_05889_));
 sky130_fd_sc_hd__nand3_1 _28428_ (.A(_05883_),
    .B(_05880_),
    .C(_05878_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_1 _28429_ (.A(_05615_),
    .B(_05617_),
    .Y(_05891_));
 sky130_fd_sc_hd__a32oi_1 _28430_ (.A1(_05738_),
    .A2(_05736_),
    .A3(_05737_),
    .B1(_05891_),
    .B2(_05607_),
    .Y(_05892_));
 sky130_fd_sc_hd__o2bb2ai_1 _28431_ (.A1_N(_05880_),
    .A2_N(_05878_),
    .B1(_05882_),
    .B2(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__nand2_1 _28432_ (.A(_05890_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__nand3_4 _28433_ (.A(_05888_),
    .B(_05889_),
    .C(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__nand2_1 _28434_ (.A(_05887_),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__nor2_2 _28435_ (.A(_05741_),
    .B(_05625_),
    .Y(_05897_));
 sky130_fd_sc_hd__a31oi_4 _28436_ (.A1(_05720_),
    .A2(_05744_),
    .A3(_05746_),
    .B1(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__nand2_4 _28437_ (.A(_05896_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__o22ai_4 _28438_ (.A1(_05625_),
    .A2(_05741_),
    .B1(_05753_),
    .B2(_05754_),
    .Y(_05900_));
 sky130_fd_sc_hd__nand3_4 _28439_ (.A(_05900_),
    .B(_05895_),
    .C(_05887_),
    .Y(_05901_));
 sky130_fd_sc_hd__nor2_4 _28440_ (.A(net448),
    .B(_05127_),
    .Y(_05902_));
 sky130_fd_sc_hd__nand2_2 _28441_ (.A(_19905_),
    .B(_05417_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand2_2 _28442_ (.A(_19901_),
    .B(_04838_),
    .Y(_05904_));
 sky130_fd_sc_hd__nor2_2 _28443_ (.A(_05903_),
    .B(_05904_),
    .Y(_05905_));
 sky130_vsdinv _28444_ (.A(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_1 _28445_ (.A(_05903_),
    .B(_05904_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_1 _28446_ (.A(_05906_),
    .B(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__nor2_2 _28447_ (.A(_05902_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__and2_1 _28448_ (.A(_05908_),
    .B(_05902_),
    .X(_05910_));
 sky130_fd_sc_hd__nor2_1 _28449_ (.A(_05909_),
    .B(_05910_),
    .Y(_05911_));
 sky130_vsdinv _28450_ (.A(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__a21o_1 _28451_ (.A1(_05899_),
    .A2(_05901_),
    .B1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__nand3_4 _28452_ (.A(_05899_),
    .B(_05901_),
    .C(_05912_),
    .Y(_05914_));
 sky130_fd_sc_hd__nand3_4 _28453_ (.A(_05913_),
    .B(_05779_),
    .C(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__nand2_1 _28454_ (.A(_05758_),
    .B(_05760_),
    .Y(_05916_));
 sky130_fd_sc_hd__a21oi_2 _28455_ (.A1(_05899_),
    .A2(_05901_),
    .B1(_05912_),
    .Y(_05917_));
 sky130_fd_sc_hd__o211a_4 _28456_ (.A1(_05910_),
    .A2(_05909_),
    .B1(_05901_),
    .C1(_05899_),
    .X(_05918_));
 sky130_fd_sc_hd__o22ai_4 _28457_ (.A1(_05762_),
    .A2(_05916_),
    .B1(_05917_),
    .B2(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__and2_4 _28458_ (.A(_05746_),
    .B(_05716_),
    .X(_05920_));
 sky130_fd_sc_hd__nor2_8 _28459_ (.A(_05920_),
    .B(_05760_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_1 _28460_ (.A(_05760_),
    .B(_05920_),
    .Y(_05922_));
 sky130_vsdinv _28461_ (.A(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__o2bb2ai_4 _28462_ (.A1_N(_05915_),
    .A2_N(_05919_),
    .B1(_05921_),
    .B2(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__nor2_4 _28463_ (.A(_05921_),
    .B(_05923_),
    .Y(_05925_));
 sky130_fd_sc_hd__nand3_4 _28464_ (.A(_05919_),
    .B(_05915_),
    .C(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__o21ai_4 _28465_ (.A1(_05784_),
    .A2(_05765_),
    .B1(_05781_),
    .Y(_05927_));
 sky130_fd_sc_hd__a21oi_2 _28466_ (.A1(_05924_),
    .A2(_05926_),
    .B1(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__a21oi_2 _28467_ (.A1(_05913_),
    .A2(_05914_),
    .B1(_05779_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_1 _28468_ (.A(_05915_),
    .B(_05925_),
    .Y(_05930_));
 sky130_fd_sc_hd__o211a_1 _28469_ (.A1(_05929_),
    .A2(_05930_),
    .B1(_05927_),
    .C1(_05924_),
    .X(_05931_));
 sky130_fd_sc_hd__o21ai_1 _28470_ (.A1(_05928_),
    .A2(_05931_),
    .B1(_05774_),
    .Y(_05932_));
 sky130_fd_sc_hd__a21o_1 _28471_ (.A1(_05924_),
    .A2(_05926_),
    .B1(_05927_),
    .X(_05933_));
 sky130_fd_sc_hd__nand3_4 _28472_ (.A(_05924_),
    .B(_05926_),
    .C(_05927_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand3_1 _28473_ (.A(_05933_),
    .B(_05783_),
    .C(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__nand3_1 _28474_ (.A(_05932_),
    .B(_05791_),
    .C(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__o22ai_2 _28475_ (.A1(_05638_),
    .A2(_05771_),
    .B1(_05928_),
    .B2(_05931_),
    .Y(_05937_));
 sky130_vsdinv _28476_ (.A(_05791_),
    .Y(_05938_));
 sky130_fd_sc_hd__nand2_2 _28477_ (.A(_05933_),
    .B(_05774_),
    .Y(_05939_));
 sky130_fd_sc_hd__nand3_1 _28478_ (.A(_05937_),
    .B(_05938_),
    .C(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_2 _28479_ (.A(_05936_),
    .B(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__a22oi_4 _28480_ (.A1(_05655_),
    .A2(_05786_),
    .B1(_05796_),
    .B2(_05793_),
    .Y(_05942_));
 sky130_fd_sc_hd__xor2_1 _28481_ (.A(_05941_),
    .B(_05942_),
    .X(_02630_));
 sky130_fd_sc_hd__or2_2 _28482_ (.A(_05612_),
    .B(_05741_),
    .X(_05943_));
 sky130_fd_sc_hd__o21ai_4 _28483_ (.A1(_05881_),
    .A2(_05943_),
    .B1(_05887_),
    .Y(_05944_));
 sky130_fd_sc_hd__a22oi_4 _28484_ (.A1(net468),
    .A2(_05283_),
    .B1(_05499_),
    .B2(_20162_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand2_4 _28485_ (.A(_20161_),
    .B(_05243_),
    .Y(_05946_));
 sky130_fd_sc_hd__nor2_8 _28486_ (.A(_05860_),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_1 _28487_ (.A(_05945_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__nand2_2 _28488_ (.A(_05506_),
    .B(_05474_),
    .Y(_05949_));
 sky130_vsdinv _28489_ (.A(_05949_),
    .Y(_05950_));
 sky130_fd_sc_hd__nand2_1 _28490_ (.A(_05948_),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__buf_6 _28491_ (.A(_19908_),
    .X(_05952_));
 sky130_fd_sc_hd__buf_8 _28492_ (.A(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__a31o_1 _28493_ (.A1(_05907_),
    .A2(_05953_),
    .A3(_05144_),
    .B1(_05905_),
    .X(_05954_));
 sky130_fd_sc_hd__o21ai_1 _28494_ (.A1(_05945_),
    .A2(_05947_),
    .B1(_05949_),
    .Y(_05955_));
 sky130_fd_sc_hd__nand3_2 _28495_ (.A(_05951_),
    .B(_05954_),
    .C(_05955_),
    .Y(_05956_));
 sky130_fd_sc_hd__nand2_1 _28496_ (.A(_05948_),
    .B(_05949_),
    .Y(_05957_));
 sky130_fd_sc_hd__a21oi_2 _28497_ (.A1(_05902_),
    .A2(_05907_),
    .B1(_05905_),
    .Y(_05958_));
 sky130_fd_sc_hd__o21ai_2 _28498_ (.A1(_05945_),
    .A2(_05947_),
    .B1(_05950_),
    .Y(_05959_));
 sky130_fd_sc_hd__nand3_4 _28499_ (.A(_05957_),
    .B(_05958_),
    .C(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__a21o_2 _28500_ (.A1(_05871_),
    .A2(_05870_),
    .B1(_05864_),
    .X(_05961_));
 sky130_fd_sc_hd__and3_1 _28501_ (.A(_05956_),
    .B(_05960_),
    .C(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_2 _28502_ (.A(_05956_),
    .X(_05963_));
 sky130_fd_sc_hd__a21o_1 _28503_ (.A1(_05960_),
    .A2(_05963_),
    .B1(_05961_),
    .X(_05964_));
 sky130_fd_sc_hd__nand2_1 _28504_ (.A(_05876_),
    .B(_05879_),
    .Y(_05965_));
 sky130_fd_sc_hd__nand2_4 _28505_ (.A(_05965_),
    .B(_05873_),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2_1 _28506_ (.A(_05964_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__nor2_2 _28507_ (.A(_05739_),
    .B(_05881_),
    .Y(_05968_));
 sky130_fd_sc_hd__a21oi_1 _28508_ (.A1(_05963_),
    .A2(_05960_),
    .B1(_05961_),
    .Y(_05969_));
 sky130_fd_sc_hd__o21bai_2 _28509_ (.A1(_05969_),
    .A2(_05962_),
    .B1_N(_05966_),
    .Y(_05970_));
 sky130_fd_sc_hd__o211ai_4 _28510_ (.A1(_05962_),
    .A2(_05967_),
    .B1(_05968_),
    .C1(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__nand3_1 _28511_ (.A(_05963_),
    .B(_05960_),
    .C(_05961_),
    .Y(_05972_));
 sky130_fd_sc_hd__a21oi_2 _28512_ (.A1(_05964_),
    .A2(_05972_),
    .B1(_05966_),
    .Y(_05973_));
 sky130_vsdinv _28513_ (.A(_05963_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand2_1 _28514_ (.A(_05960_),
    .B(_05961_),
    .Y(_05975_));
 sky130_fd_sc_hd__o211a_1 _28515_ (.A1(_05974_),
    .A2(_05975_),
    .B1(_05966_),
    .C1(_05964_),
    .X(_05976_));
 sky130_fd_sc_hd__o22ai_4 _28516_ (.A1(_05739_),
    .A2(_05881_),
    .B1(_05973_),
    .B2(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__clkbuf_2 _28517_ (.A(_05377_),
    .X(_05978_));
 sky130_fd_sc_hd__buf_6 _28518_ (.A(_05571_),
    .X(_05979_));
 sky130_fd_sc_hd__a22oi_4 _28519_ (.A1(_05816_),
    .A2(_05693_),
    .B1(net447),
    .B2(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__buf_6 _28520_ (.A(_05372_),
    .X(_05981_));
 sky130_fd_sc_hd__and4_4 _28521_ (.A(_05213_),
    .B(_05558_),
    .C(_05698_),
    .D(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__a211o_1 _28522_ (.A1(_19938_),
    .A2(_20139_),
    .B1(_05980_),
    .C1(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__a21oi_4 _28523_ (.A1(_05807_),
    .A2(_05802_),
    .B1(_05800_),
    .Y(_05984_));
 sky130_fd_sc_hd__buf_6 _28524_ (.A(\pcpi_mul.rs1[12] ),
    .X(_05985_));
 sky130_fd_sc_hd__buf_6 _28525_ (.A(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__nand2_2 _28526_ (.A(_05192_),
    .B(_05986_),
    .Y(_05987_));
 sky130_vsdinv _28527_ (.A(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__o21ai_2 _28528_ (.A1(_05980_),
    .A2(_05982_),
    .B1(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__nand3_4 _28529_ (.A(_05983_),
    .B(_05984_),
    .C(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__buf_6 _28530_ (.A(_05571_),
    .X(_05991_));
 sky130_fd_sc_hd__a22o_2 _28531_ (.A1(_05816_),
    .A2(_05693_),
    .B1(_05674_),
    .B2(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__nand3b_4 _28532_ (.A_N(_05982_),
    .B(_05988_),
    .C(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__o21ai_4 _28533_ (.A1(_05801_),
    .A2(_05798_),
    .B1(_05806_),
    .Y(_05994_));
 sky130_fd_sc_hd__o21ai_4 _28534_ (.A1(_05980_),
    .A2(_05982_),
    .B1(_05987_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand3_4 _28535_ (.A(_05993_),
    .B(_05994_),
    .C(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__nand2_1 _28536_ (.A(_05990_),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__buf_6 _28537_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05998_));
 sky130_fd_sc_hd__clkbuf_8 _28538_ (.A(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__and4_2 _28539_ (.A(_05240_),
    .B(_05284_),
    .C(_05999_),
    .D(_05835_),
    .X(_06000_));
 sky130_fd_sc_hd__nand2_1 _28540_ (.A(_05174_),
    .B(_05823_),
    .Y(_06001_));
 sky130_fd_sc_hd__o21a_1 _28541_ (.A1(_05250_),
    .A2(_05813_),
    .B1(_06001_),
    .X(_06002_));
 sky130_vsdinv _28542_ (.A(\pcpi_mul.rs1[9] ),
    .Y(_06003_));
 sky130_fd_sc_hd__buf_8 _28543_ (.A(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__nor2_1 _28544_ (.A(_05186_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__o21bai_1 _28545_ (.A1(_06000_),
    .A2(_06002_),
    .B1_N(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__o21ai_1 _28546_ (.A1(_05151_),
    .A2(_05813_),
    .B1(_06001_),
    .Y(_06007_));
 sky130_fd_sc_hd__nand3b_2 _28547_ (.A_N(_06000_),
    .B(_06005_),
    .C(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_2 _28548_ (.A(_06006_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2_2 _28549_ (.A(_05997_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2_2 _28550_ (.A(_05819_),
    .B(_05838_),
    .Y(_06011_));
 sky130_fd_sc_hd__and2_1 _28551_ (.A(_06011_),
    .B(_05811_),
    .X(_06012_));
 sky130_fd_sc_hd__and2_1 _28552_ (.A(_06006_),
    .B(_06008_),
    .X(_06013_));
 sky130_fd_sc_hd__nand3_4 _28553_ (.A(_06013_),
    .B(_05990_),
    .C(_05996_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand3_4 _28554_ (.A(_06010_),
    .B(_06012_),
    .C(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_1 _28555_ (.A(_05997_),
    .B(_06013_),
    .Y(_06016_));
 sky130_fd_sc_hd__nand2_1 _28556_ (.A(_06011_),
    .B(_05811_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand3_2 _28557_ (.A(_05990_),
    .B(_06009_),
    .C(_05996_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand3_4 _28558_ (.A(_06016_),
    .B(_06017_),
    .C(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__nor2_8 _28559_ (.A(_05829_),
    .B(_05848_),
    .Y(_06020_));
 sky130_fd_sc_hd__a21oi_1 _28560_ (.A1(_06015_),
    .A2(_06019_),
    .B1(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand3_4 _28561_ (.A(_06015_),
    .B(_06019_),
    .C(_06020_),
    .Y(_06022_));
 sky130_vsdinv _28562_ (.A(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__o2bb2ai_1 _28563_ (.A1_N(_05971_),
    .A2_N(_05977_),
    .B1(_06021_),
    .B2(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__clkbuf_4 _28564_ (.A(_05976_),
    .X(_06025_));
 sky130_fd_sc_hd__nand2_1 _28565_ (.A(_05970_),
    .B(_05968_),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2_1 _28566_ (.A(_06015_),
    .B(_06019_),
    .Y(_06027_));
 sky130_vsdinv _28567_ (.A(_06020_),
    .Y(_06028_));
 sky130_fd_sc_hd__nand2_1 _28568_ (.A(_06027_),
    .B(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__o2111ai_4 _28569_ (.A1(_06025_),
    .A2(_06026_),
    .B1(_06029_),
    .C1(_06022_),
    .D1(_05977_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand3b_4 _28570_ (.A_N(_05944_),
    .B(_06024_),
    .C(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__a21oi_1 _28571_ (.A1(_06015_),
    .A2(_06019_),
    .B1(_06028_),
    .Y(_06032_));
 sky130_fd_sc_hd__nor2_1 _28572_ (.A(_06020_),
    .B(_06027_),
    .Y(_06033_));
 sky130_fd_sc_hd__o2bb2ai_2 _28573_ (.A1_N(_05971_),
    .A2_N(_05977_),
    .B1(_06032_),
    .B2(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__and3_1 _28574_ (.A(_06010_),
    .B(_06012_),
    .C(_06014_),
    .X(_06035_));
 sky130_fd_sc_hd__nand2_2 _28575_ (.A(_06019_),
    .B(_06028_),
    .Y(_06036_));
 sky130_fd_sc_hd__nand2_1 _28576_ (.A(_06027_),
    .B(_06020_),
    .Y(_06037_));
 sky130_fd_sc_hd__o2111ai_4 _28577_ (.A1(_06035_),
    .A2(_06036_),
    .B1(_05971_),
    .C1(_06037_),
    .D1(_05977_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand3_4 _28578_ (.A(_06034_),
    .B(_06038_),
    .C(_05944_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_2 _28579_ (.A(net455),
    .B(_20178_),
    .Y(_06040_));
 sky130_fd_sc_hd__clkbuf_4 _28580_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06041_));
 sky130_fd_sc_hd__buf_4 _28581_ (.A(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__nand2_1 _28582_ (.A(_06042_),
    .B(_20174_),
    .Y(_06043_));
 sky130_fd_sc_hd__buf_4 _28583_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06044_));
 sky130_fd_sc_hd__buf_6 _28584_ (.A(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__buf_8 _28585_ (.A(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__nand3b_4 _28586_ (.A_N(_06043_),
    .B(_06046_),
    .C(_20172_),
    .Y(_06047_));
 sky130_fd_sc_hd__buf_6 _28587_ (.A(_19901_),
    .X(_06048_));
 sky130_fd_sc_hd__buf_8 _28588_ (.A(_19905_),
    .X(_06049_));
 sky130_fd_sc_hd__a22o_1 _28589_ (.A1(_06048_),
    .A2(_05418_),
    .B1(_06049_),
    .B2(_05181_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_4 _28590_ (.A(\pcpi_mul.rs2[9] ),
    .X(_06051_));
 sky130_fd_sc_hd__buf_8 _28591_ (.A(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__nand2_1 _28592_ (.A(_06052_),
    .B(_05177_),
    .Y(_06053_));
 sky130_vsdinv _28593_ (.A(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a21oi_4 _28594_ (.A1(_06047_),
    .A2(_06050_),
    .B1(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__and3_1 _28595_ (.A(_06047_),
    .B(_06054_),
    .C(_06050_),
    .X(_06056_));
 sky130_fd_sc_hd__nor3_4 _28596_ (.A(_06040_),
    .B(_06055_),
    .C(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__o21a_4 _28597_ (.A1(_06055_),
    .A2(_06056_),
    .B1(_06040_),
    .X(_06058_));
 sky130_fd_sc_hd__nor2_8 _28598_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__a21o_1 _28599_ (.A1(_06031_),
    .A2(_06039_),
    .B1(_06059_),
    .X(_06060_));
 sky130_fd_sc_hd__nand3_4 _28600_ (.A(_06031_),
    .B(_06039_),
    .C(_06059_),
    .Y(_06061_));
 sky130_fd_sc_hd__a21oi_4 _28601_ (.A1(_06060_),
    .A2(_06061_),
    .B1(_05918_),
    .Y(_06062_));
 sky130_fd_sc_hd__a21oi_4 _28602_ (.A1(_06031_),
    .A2(_06039_),
    .B1(_06059_),
    .Y(_06063_));
 sky130_vsdinv _28603_ (.A(_06061_),
    .Y(_06064_));
 sky130_fd_sc_hd__nor3_4 _28604_ (.A(_05914_),
    .B(_06063_),
    .C(_06064_),
    .Y(_06065_));
 sky130_vsdinv _28605_ (.A(_05852_),
    .Y(_06066_));
 sky130_fd_sc_hd__a21oi_4 _28606_ (.A1(_05856_),
    .A2(_05843_),
    .B1(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__nor2_4 _28607_ (.A(_06067_),
    .B(_05901_),
    .Y(_06068_));
 sky130_fd_sc_hd__and2_1 _28608_ (.A(_05901_),
    .B(_06067_),
    .X(_06069_));
 sky130_fd_sc_hd__or2_2 _28609_ (.A(_06068_),
    .B(_06069_),
    .X(_06070_));
 sky130_vsdinv _28610_ (.A(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__o21ai_2 _28611_ (.A1(_06062_),
    .A2(_06065_),
    .B1(_06071_),
    .Y(_06072_));
 sky130_vsdinv _28612_ (.A(_05925_),
    .Y(_06073_));
 sky130_fd_sc_hd__o21a_1 _28613_ (.A1(_05929_),
    .A2(_06073_),
    .B1(_05915_),
    .X(_06074_));
 sky130_fd_sc_hd__o21ai_1 _28614_ (.A1(_06063_),
    .A2(_06064_),
    .B1(_05914_),
    .Y(_06075_));
 sky130_fd_sc_hd__nand3_4 _28615_ (.A(_06060_),
    .B(_05918_),
    .C(_06061_),
    .Y(_06076_));
 sky130_fd_sc_hd__nand3_2 _28616_ (.A(_06075_),
    .B(_06070_),
    .C(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand3_4 _28617_ (.A(_06072_),
    .B(_06074_),
    .C(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2_4 _28618_ (.A(_06078_),
    .B(_05921_),
    .Y(_06079_));
 sky130_fd_sc_hd__o22ai_2 _28619_ (.A1(_06068_),
    .A2(_06069_),
    .B1(_06062_),
    .B2(_06065_),
    .Y(_06080_));
 sky130_fd_sc_hd__nand3_1 _28620_ (.A(_06071_),
    .B(_06075_),
    .C(_06076_),
    .Y(_06081_));
 sky130_fd_sc_hd__o21ai_1 _28621_ (.A1(_05929_),
    .A2(_06073_),
    .B1(_05915_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand3_2 _28622_ (.A(_06080_),
    .B(_06081_),
    .C(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2_1 _28623_ (.A(_06078_),
    .B(_06083_),
    .Y(_06084_));
 sky130_vsdinv _28624_ (.A(_05921_),
    .Y(_06085_));
 sky130_fd_sc_hd__a22oi_4 _28625_ (.A1(_05939_),
    .A2(_05934_),
    .B1(_06084_),
    .B2(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__o2bb2ai_1 _28626_ (.A1_N(_06083_),
    .A2_N(_06078_),
    .B1(_05760_),
    .B2(_05920_),
    .Y(_06087_));
 sky130_fd_sc_hd__nand2_1 _28627_ (.A(_05939_),
    .B(_05934_),
    .Y(_06088_));
 sky130_fd_sc_hd__a21oi_2 _28628_ (.A1(_06087_),
    .A2(_06079_),
    .B1(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__a21oi_4 _28629_ (.A1(_06079_),
    .A2(_06086_),
    .B1(_06089_),
    .Y(_06090_));
 sky130_vsdinv _28630_ (.A(_05939_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand2_1 _28631_ (.A(_05937_),
    .B(_05938_),
    .Y(_06092_));
 sky130_fd_sc_hd__o22ai_4 _28632_ (.A1(_06091_),
    .A2(_06092_),
    .B1(_05941_),
    .B2(_05942_),
    .Y(_06093_));
 sky130_fd_sc_hd__xor2_1 _28633_ (.A(_06090_),
    .B(_06093_),
    .X(_02631_));
 sky130_fd_sc_hd__nand2_2 _28634_ (.A(_06038_),
    .B(_05971_),
    .Y(_06094_));
 sky130_fd_sc_hd__buf_8 _28635_ (.A(_05501_),
    .X(_06095_));
 sky130_fd_sc_hd__buf_8 _28636_ (.A(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__buf_4 _28637_ (.A(_05412_),
    .X(_06097_));
 sky130_fd_sc_hd__buf_8 _28638_ (.A(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__a22oi_4 _28639_ (.A1(_06096_),
    .A2(_20163_),
    .B1(_06098_),
    .B2(_20159_),
    .Y(_06099_));
 sky130_fd_sc_hd__clkbuf_8 _28640_ (.A(_05722_),
    .X(_06100_));
 sky130_fd_sc_hd__nand3_4 _28641_ (.A(_06100_),
    .B(_19915_),
    .C(_05481_),
    .Y(_06101_));
 sky130_fd_sc_hd__nor2_4 _28642_ (.A(_05580_),
    .B(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand2_2 _28643_ (.A(_05866_),
    .B(_05573_),
    .Y(_06103_));
 sky130_vsdinv _28644_ (.A(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__o21ai_2 _28645_ (.A1(_06099_),
    .A2(_06102_),
    .B1(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__buf_2 _28646_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_8 _28647_ (.A(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__and4_1 _28648_ (.A(_19902_),
    .B(_06107_),
    .C(_05181_),
    .D(_05418_),
    .X(_06108_));
 sky130_fd_sc_hd__a21oi_2 _28649_ (.A1(_06050_),
    .A2(_06054_),
    .B1(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__buf_6 _28650_ (.A(_05412_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_8 _28651_ (.A(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__a22o_2 _28652_ (.A1(_05858_),
    .A2(_20163_),
    .B1(_06111_),
    .B2(_20159_),
    .X(_06112_));
 sky130_fd_sc_hd__o211ai_2 _28653_ (.A1(_05296_),
    .A2(_06101_),
    .B1(_06103_),
    .C1(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand3_4 _28654_ (.A(_06105_),
    .B(_06109_),
    .C(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__o21ai_2 _28655_ (.A1(_06099_),
    .A2(_06102_),
    .B1(_06103_),
    .Y(_06115_));
 sky130_fd_sc_hd__o211ai_2 _28656_ (.A1(_05296_),
    .A2(_06101_),
    .B1(_06104_),
    .C1(_06112_),
    .Y(_06116_));
 sky130_fd_sc_hd__buf_4 _28657_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06117_));
 sky130_fd_sc_hd__buf_6 _28658_ (.A(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__buf_6 _28659_ (.A(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__a22oi_2 _28660_ (.A1(_06119_),
    .A2(_05147_),
    .B1(_06046_),
    .B2(_20172_),
    .Y(_06120_));
 sky130_fd_sc_hd__o21ai_2 _28661_ (.A1(_06053_),
    .A2(_06120_),
    .B1(_06047_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand3_4 _28662_ (.A(_06115_),
    .B(_06116_),
    .C(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__nand2_1 _28663_ (.A(_06114_),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__nor2_2 _28664_ (.A(_05949_),
    .B(_05945_),
    .Y(_06124_));
 sky130_fd_sc_hd__nor2_4 _28665_ (.A(_05947_),
    .B(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_4 _28666_ (.A(_06123_),
    .B(_06125_),
    .Y(_06126_));
 sky130_vsdinv _28667_ (.A(_06125_),
    .Y(_06127_));
 sky130_fd_sc_hd__nand3_4 _28668_ (.A(_06127_),
    .B(_06114_),
    .C(_06122_),
    .Y(_06128_));
 sky130_fd_sc_hd__a21oi_4 _28669_ (.A1(_06126_),
    .A2(_06128_),
    .B1(_06057_),
    .Y(_06129_));
 sky130_fd_sc_hd__and3_1 _28670_ (.A(_06126_),
    .B(_06057_),
    .C(_06128_),
    .X(_06130_));
 sky130_fd_sc_hd__and2_2 _28671_ (.A(_05975_),
    .B(_05963_),
    .X(_06131_));
 sky130_fd_sc_hd__o21ai_4 _28672_ (.A1(_06129_),
    .A2(_06130_),
    .B1(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__a21o_1 _28673_ (.A1(_06126_),
    .A2(_06128_),
    .B1(_06057_),
    .X(_06133_));
 sky130_fd_sc_hd__nand3_4 _28674_ (.A(_06126_),
    .B(_06057_),
    .C(_06128_),
    .Y(_06134_));
 sky130_fd_sc_hd__nand2_1 _28675_ (.A(_05975_),
    .B(_05963_),
    .Y(_06135_));
 sky130_fd_sc_hd__nand3_4 _28676_ (.A(_06133_),
    .B(_06134_),
    .C(_06135_),
    .Y(_06136_));
 sky130_fd_sc_hd__a21oi_4 _28677_ (.A1(_06132_),
    .A2(_06136_),
    .B1(_06025_),
    .Y(_06137_));
 sky130_fd_sc_hd__and3_1 _28678_ (.A(_06132_),
    .B(_06025_),
    .C(_06136_),
    .X(_06138_));
 sky130_fd_sc_hd__a22oi_4 _28679_ (.A1(_05229_),
    .A2(_05832_),
    .B1(_05805_),
    .B2(net454),
    .Y(_06139_));
 sky130_fd_sc_hd__nand3_4 _28680_ (.A(_19920_),
    .B(_05298_),
    .C(_20152_),
    .Y(_06140_));
 sky130_fd_sc_hd__nor2_8 _28681_ (.A(_06004_),
    .B(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__buf_4 _28682_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06142_));
 sky130_fd_sc_hd__buf_8 _28683_ (.A(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__nand2_4 _28684_ (.A(_05192_),
    .B(_06143_),
    .Y(_06144_));
 sky130_vsdinv _28685_ (.A(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__o21ai_2 _28686_ (.A1(_06139_),
    .A2(_06141_),
    .B1(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__a21oi_4 _28687_ (.A1(_05992_),
    .A2(_05988_),
    .B1(_05982_),
    .Y(_06147_));
 sky130_fd_sc_hd__clkbuf_4 _28688_ (.A(_05555_),
    .X(_06148_));
 sky130_fd_sc_hd__a22o_2 _28689_ (.A1(_05229_),
    .A2(_05979_),
    .B1(net447),
    .B2(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__o211ai_4 _28690_ (.A1(_06004_),
    .A2(_06140_),
    .B1(_06144_),
    .C1(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__buf_6 _28691_ (.A(_05985_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_4 _28692_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06152_));
 sky130_fd_sc_hd__buf_6 _28693_ (.A(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__buf_6 _28694_ (.A(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_8 _28695_ (.A(_06151_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__nor2_4 _28696_ (.A(_05130_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__nand2_2 _28697_ (.A(_19929_),
    .B(_20147_),
    .Y(_06157_));
 sky130_fd_sc_hd__a22o_2 _28698_ (.A1(_05140_),
    .A2(_20143_),
    .B1(_19935_),
    .B2(_20139_),
    .X(_06158_));
 sky130_fd_sc_hd__nand3b_4 _28699_ (.A_N(_06156_),
    .B(_06157_),
    .C(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__o21ai_4 _28700_ (.A1(_05130_),
    .A2(_06155_),
    .B1(_06158_),
    .Y(_06160_));
 sky130_fd_sc_hd__nand3_4 _28701_ (.A(_06160_),
    .B(_19929_),
    .C(_20147_),
    .Y(_06161_));
 sky130_fd_sc_hd__a32oi_4 _28702_ (.A1(_06146_),
    .A2(_06147_),
    .A3(_06150_),
    .B1(_06159_),
    .B2(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__nand2_1 _28703_ (.A(_06149_),
    .B(_06145_),
    .Y(_06163_));
 sky130_fd_sc_hd__o21ai_2 _28704_ (.A1(_06139_),
    .A2(_06141_),
    .B1(_06144_),
    .Y(_06164_));
 sky130_fd_sc_hd__a21o_1 _28705_ (.A1(_05992_),
    .A2(_05988_),
    .B1(_05982_),
    .X(_06165_));
 sky130_fd_sc_hd__o211ai_4 _28706_ (.A1(_06141_),
    .A2(_06163_),
    .B1(_06164_),
    .C1(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_2 _28707_ (.A(_06162_),
    .B(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__nand3_1 _28708_ (.A(_06146_),
    .B(_06147_),
    .C(_06150_),
    .Y(_06168_));
 sky130_fd_sc_hd__nand2_1 _28709_ (.A(_06161_),
    .B(_06159_),
    .Y(_06169_));
 sky130_fd_sc_hd__a21o_1 _28710_ (.A1(_06166_),
    .A2(_06168_),
    .B1(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__a21oi_4 _28711_ (.A1(_05993_),
    .A2(_05995_),
    .B1(_05994_),
    .Y(_06171_));
 sky130_fd_sc_hd__o21ai_4 _28712_ (.A1(_06009_),
    .A2(_06171_),
    .B1(_05996_),
    .Y(_06172_));
 sky130_fd_sc_hd__a21oi_1 _28713_ (.A1(_06167_),
    .A2(_06170_),
    .B1(_06172_),
    .Y(_06173_));
 sky130_vsdinv _28714_ (.A(_06166_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand2_1 _28715_ (.A(_06169_),
    .B(_06168_),
    .Y(_06175_));
 sky130_fd_sc_hd__o211a_1 _28716_ (.A1(_06174_),
    .A2(_06175_),
    .B1(_06170_),
    .C1(_06172_),
    .X(_06176_));
 sky130_vsdinv _28717_ (.A(_06008_),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_2 _28718_ (.A(_06000_),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__o21ai_2 _28719_ (.A1(_06173_),
    .A2(_06176_),
    .B1(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__a21o_1 _28720_ (.A1(_06167_),
    .A2(_06170_),
    .B1(_06172_),
    .X(_06180_));
 sky130_vsdinv _28721_ (.A(_06178_),
    .Y(_06181_));
 sky130_fd_sc_hd__nand3_4 _28722_ (.A(_06167_),
    .B(_06172_),
    .C(_06170_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand3_4 _28723_ (.A(_06180_),
    .B(_06181_),
    .C(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__and2_1 _28724_ (.A(_06179_),
    .B(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__o21ai_2 _28725_ (.A1(_06137_),
    .A2(_06138_),
    .B1(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__a21o_1 _28726_ (.A1(_06132_),
    .A2(_06136_),
    .B1(_06025_),
    .X(_06186_));
 sky130_fd_sc_hd__nand2_4 _28727_ (.A(_06179_),
    .B(_06183_),
    .Y(_06187_));
 sky130_fd_sc_hd__nand3_4 _28728_ (.A(_06132_),
    .B(_06025_),
    .C(_06136_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand3_2 _28729_ (.A(_06186_),
    .B(_06187_),
    .C(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand3b_4 _28730_ (.A_N(_06094_),
    .B(_06185_),
    .C(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__o21ai_2 _28731_ (.A1(_06137_),
    .A2(_06138_),
    .B1(_06187_),
    .Y(_06191_));
 sky130_fd_sc_hd__nand3_2 _28732_ (.A(_06184_),
    .B(_06186_),
    .C(_06188_),
    .Y(_06192_));
 sky130_fd_sc_hd__nand3_4 _28733_ (.A(_06191_),
    .B(_06192_),
    .C(_06094_),
    .Y(_06193_));
 sky130_fd_sc_hd__nand2_2 _28734_ (.A(_06190_),
    .B(_06193_),
    .Y(_06194_));
 sky130_fd_sc_hd__a22oi_4 _28735_ (.A1(_06048_),
    .A2(_05181_),
    .B1(_06049_),
    .B2(_20169_),
    .Y(_06195_));
 sky130_fd_sc_hd__buf_8 _28736_ (.A(_06044_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_4 _28737_ (.A(_05178_),
    .X(_06197_));
 sky130_fd_sc_hd__and4_1 _28738_ (.A(_06042_),
    .B(_06196_),
    .C(_05177_),
    .D(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__buf_8 _28739_ (.A(_20164_),
    .X(_06199_));
 sky130_fd_sc_hd__nand2_2 _28740_ (.A(_19909_),
    .B(_06199_),
    .Y(_06200_));
 sky130_vsdinv _28741_ (.A(_06200_),
    .Y(_06201_));
 sky130_fd_sc_hd__o21ai_2 _28742_ (.A1(_06195_),
    .A2(_06198_),
    .B1(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__nand2_1 _28743_ (.A(_06042_),
    .B(_06197_),
    .Y(_06203_));
 sky130_fd_sc_hd__nand3b_4 _28744_ (.A_N(_06203_),
    .B(_06046_),
    .C(_20169_),
    .Y(_06204_));
 sky130_fd_sc_hd__a22o_2 _28745_ (.A1(_19902_),
    .A2(_05179_),
    .B1(_19906_),
    .B2(_05183_),
    .X(_06205_));
 sky130_fd_sc_hd__nand3_4 _28746_ (.A(_06204_),
    .B(_06205_),
    .C(_06200_),
    .Y(_06206_));
 sky130_fd_sc_hd__buf_6 _28747_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_8 _28748_ (.A(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__nand2_1 _28749_ (.A(_06208_),
    .B(_05230_),
    .Y(_06209_));
 sky130_fd_sc_hd__nand2_1 _28750_ (.A(_19899_),
    .B(_20174_),
    .Y(_06210_));
 sky130_fd_sc_hd__or2_2 _28751_ (.A(_06209_),
    .B(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__nand2_1 _28752_ (.A(_06209_),
    .B(_06210_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_2 _28753_ (.A(_06211_),
    .B(_06212_),
    .Y(_06213_));
 sky130_fd_sc_hd__a21oi_4 _28754_ (.A1(_06202_),
    .A2(_06206_),
    .B1(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__and3_1 _28755_ (.A(_06213_),
    .B(_06202_),
    .C(_06206_),
    .X(_06215_));
 sky130_fd_sc_hd__or2_4 _28756_ (.A(_06214_),
    .B(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__nand2_2 _28757_ (.A(_06194_),
    .B(_06216_),
    .Y(_06217_));
 sky130_vsdinv _28758_ (.A(_06216_),
    .Y(_06218_));
 sky130_fd_sc_hd__nand3_4 _28759_ (.A(_06190_),
    .B(_06193_),
    .C(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__nand3_4 _28760_ (.A(_06217_),
    .B(_06064_),
    .C(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__a21o_1 _28761_ (.A1(_06217_),
    .A2(_06219_),
    .B1(_06064_),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _28762_ (.A(_06036_),
    .B(_06015_),
    .Y(_06222_));
 sky130_fd_sc_hd__and2_1 _28763_ (.A(_06039_),
    .B(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__nor2_1 _28764_ (.A(_06222_),
    .B(_06039_),
    .Y(_06224_));
 sky130_fd_sc_hd__o2bb2ai_1 _28765_ (.A1_N(_06220_),
    .A2_N(_06221_),
    .B1(_06223_),
    .B2(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__o21a_1 _28766_ (.A1(_06070_),
    .A2(_06062_),
    .B1(_06076_),
    .X(_06226_));
 sky130_fd_sc_hd__nor2_2 _28767_ (.A(_06224_),
    .B(_06223_),
    .Y(_06227_));
 sky130_fd_sc_hd__nand3_1 _28768_ (.A(_06221_),
    .B(_06227_),
    .C(_06220_),
    .Y(_06228_));
 sky130_fd_sc_hd__nand3_2 _28769_ (.A(_06225_),
    .B(_06226_),
    .C(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__and2_1 _28770_ (.A(_06229_),
    .B(_06068_),
    .X(_06230_));
 sky130_fd_sc_hd__nand2_1 _28771_ (.A(_06221_),
    .B(_06220_),
    .Y(_06231_));
 sky130_fd_sc_hd__nand2_1 _28772_ (.A(_06231_),
    .B(_06227_),
    .Y(_06232_));
 sky130_vsdinv _28773_ (.A(_06226_),
    .Y(_06233_));
 sky130_vsdinv _28774_ (.A(_06227_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand3_1 _28775_ (.A(_06221_),
    .B(_06234_),
    .C(_06220_),
    .Y(_06235_));
 sky130_fd_sc_hd__nand3_2 _28776_ (.A(_06232_),
    .B(_06233_),
    .C(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__a21o_1 _28777_ (.A1(_06236_),
    .A2(_06229_),
    .B1(_06068_),
    .X(_06237_));
 sky130_fd_sc_hd__nand2_1 _28778_ (.A(_06079_),
    .B(_06083_),
    .Y(_06238_));
 sky130_fd_sc_hd__nand2_1 _28779_ (.A(_06237_),
    .B(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__a21oi_1 _28780_ (.A1(_06236_),
    .A2(_06229_),
    .B1(_06068_),
    .Y(_06240_));
 sky130_fd_sc_hd__o21bai_1 _28781_ (.A1(_06230_),
    .A2(_06240_),
    .B1_N(_06238_),
    .Y(_06241_));
 sky130_fd_sc_hd__o21ai_2 _28782_ (.A1(_06230_),
    .A2(_06239_),
    .B1(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__a22oi_4 _28783_ (.A1(_06079_),
    .A2(_06086_),
    .B1(_06093_),
    .B2(_06090_),
    .Y(_06243_));
 sky130_fd_sc_hd__xor2_1 _28784_ (.A(_06242_),
    .B(_06243_),
    .X(_02632_));
 sky130_fd_sc_hd__a21bo_1 _28785_ (.A1(_06221_),
    .A2(_06234_),
    .B1_N(_06220_),
    .X(_06244_));
 sky130_fd_sc_hd__a21oi_4 _28786_ (.A1(_06112_),
    .A2(_06104_),
    .B1(_06102_),
    .Y(_06245_));
 sky130_fd_sc_hd__a22oi_4 _28787_ (.A1(net467),
    .A2(_05675_),
    .B1(_06111_),
    .B2(_05697_),
    .Y(_06246_));
 sky130_vsdinv _28788_ (.A(_20154_),
    .Y(_06247_));
 sky130_fd_sc_hd__clkbuf_2 _28789_ (.A(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__buf_6 _28790_ (.A(_05664_),
    .X(_06249_));
 sky130_fd_sc_hd__nand3_4 _28791_ (.A(_06095_),
    .B(_05499_),
    .C(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nor2_8 _28792_ (.A(net446),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__nand2_2 _28793_ (.A(_05506_),
    .B(_05831_),
    .Y(_06252_));
 sky130_vsdinv _28794_ (.A(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__o21ai_2 _28795_ (.A1(_06246_),
    .A2(_06251_),
    .B1(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__a21oi_2 _28796_ (.A1(_06205_),
    .A2(_06201_),
    .B1(_06198_),
    .Y(_06255_));
 sky130_fd_sc_hd__buf_8 _28797_ (.A(net446),
    .X(_06256_));
 sky130_fd_sc_hd__a22o_2 _28798_ (.A1(_05858_),
    .A2(_20159_),
    .B1(_05414_),
    .B2(_05697_),
    .X(_06257_));
 sky130_fd_sc_hd__o211ai_4 _28799_ (.A1(_06256_),
    .A2(_06250_),
    .B1(_06252_),
    .C1(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__nand3_4 _28800_ (.A(_06254_),
    .B(_06255_),
    .C(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__o21ai_2 _28801_ (.A1(_06246_),
    .A2(_06251_),
    .B1(_06252_),
    .Y(_06260_));
 sky130_fd_sc_hd__o211ai_4 _28802_ (.A1(_06256_),
    .A2(_06250_),
    .B1(_06253_),
    .C1(_06257_),
    .Y(_06261_));
 sky130_fd_sc_hd__o21ai_2 _28803_ (.A1(_06200_),
    .A2(_06195_),
    .B1(_06204_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand3_4 _28804_ (.A(_06260_),
    .B(_06261_),
    .C(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__nand2_2 _28805_ (.A(_06259_),
    .B(_06263_),
    .Y(_06264_));
 sky130_vsdinv _28806_ (.A(_06245_),
    .Y(_06265_));
 sky130_fd_sc_hd__nand3_4 _28807_ (.A(_06259_),
    .B(_06263_),
    .C(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_2 _28808_ (.A(_06266_),
    .B(_06214_),
    .Y(_06267_));
 sky130_fd_sc_hd__a21oi_4 _28809_ (.A1(_06245_),
    .A2(_06264_),
    .B1(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_2 _28810_ (.A(_06264_),
    .B(_06245_),
    .Y(_06269_));
 sky130_fd_sc_hd__a21oi_4 _28811_ (.A1(_06269_),
    .A2(_06266_),
    .B1(_06214_),
    .Y(_06270_));
 sky130_fd_sc_hd__nand2_1 _28812_ (.A(_06127_),
    .B(_06114_),
    .Y(_06271_));
 sky130_fd_sc_hd__nand2_2 _28813_ (.A(_06271_),
    .B(_06122_),
    .Y(_06272_));
 sky130_fd_sc_hd__o21ai_4 _28814_ (.A1(_06268_),
    .A2(_06270_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nand2_1 _28815_ (.A(_06131_),
    .B(_06134_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand2_2 _28816_ (.A(_06274_),
    .B(_06133_),
    .Y(_06275_));
 sky130_fd_sc_hd__a21o_2 _28817_ (.A1(_06245_),
    .A2(_06264_),
    .B1(_06267_),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_1 _28818_ (.A(_06269_),
    .B(_06266_),
    .Y(_06277_));
 sky130_vsdinv _28819_ (.A(_06214_),
    .Y(_06278_));
 sky130_fd_sc_hd__nand2_2 _28820_ (.A(_06277_),
    .B(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__and2_2 _28821_ (.A(_06271_),
    .B(_06122_),
    .X(_06280_));
 sky130_fd_sc_hd__nand3_4 _28822_ (.A(_06276_),
    .B(_06279_),
    .C(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand3_4 _28823_ (.A(_06273_),
    .B(_06275_),
    .C(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__o21ai_2 _28824_ (.A1(_06268_),
    .A2(_06270_),
    .B1(_06280_),
    .Y(_06283_));
 sky130_fd_sc_hd__o21ai_2 _28825_ (.A1(_06131_),
    .A2(_06129_),
    .B1(_06134_),
    .Y(_06284_));
 sky130_fd_sc_hd__nand3_2 _28826_ (.A(_06276_),
    .B(_06279_),
    .C(_06272_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand3_4 _28827_ (.A(_06283_),
    .B(_06284_),
    .C(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__clkinv_8 _28828_ (.A(_20144_),
    .Y(_06287_));
 sky130_fd_sc_hd__clkbuf_8 _28829_ (.A(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__buf_8 _28830_ (.A(_20148_),
    .X(_06289_));
 sky130_fd_sc_hd__nand3_4 _28831_ (.A(_05797_),
    .B(_05298_),
    .C(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__a22o_4 _28832_ (.A1(_05213_),
    .A2(_05699_),
    .B1(_05558_),
    .B2(_05835_),
    .X(_06291_));
 sky130_fd_sc_hd__o21ai_1 _28833_ (.A1(_06288_),
    .A2(_06290_),
    .B1(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__clkbuf_4 _28834_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06293_));
 sky130_fd_sc_hd__buf_6 _28835_ (.A(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__nand2_2 _28836_ (.A(_05307_),
    .B(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_1 _28837_ (.A(_06292_),
    .B(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__buf_2 _28838_ (.A(_06287_),
    .X(_06297_));
 sky130_fd_sc_hd__buf_6 _28839_ (.A(net445),
    .X(_06298_));
 sky130_vsdinv _28840_ (.A(_06295_),
    .Y(_06299_));
 sky130_fd_sc_hd__o211ai_2 _28841_ (.A1(_06298_),
    .A2(_06290_),
    .B1(_06299_),
    .C1(_06291_),
    .Y(_06300_));
 sky130_fd_sc_hd__o22ai_4 _28842_ (.A1(_06004_),
    .A2(_06140_),
    .B1(_06144_),
    .B2(_06139_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand3_4 _28843_ (.A(_06296_),
    .B(_06300_),
    .C(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__nand2_2 _28844_ (.A(_06292_),
    .B(_06299_),
    .Y(_06303_));
 sky130_fd_sc_hd__a21oi_4 _28845_ (.A1(_06149_),
    .A2(_06145_),
    .B1(_06141_),
    .Y(_06304_));
 sky130_fd_sc_hd__o211ai_4 _28846_ (.A1(_06298_),
    .A2(_06290_),
    .B1(_06295_),
    .C1(_06291_),
    .Y(_06305_));
 sky130_fd_sc_hd__nand3_4 _28847_ (.A(_06303_),
    .B(_06304_),
    .C(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__buf_8 _28848_ (.A(_05812_),
    .X(_06307_));
 sky130_fd_sc_hd__buf_6 _28849_ (.A(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__buf_4 _28850_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06309_));
 sky130_fd_sc_hd__clkbuf_2 _28851_ (.A(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__buf_6 _28852_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06311_));
 sky130_fd_sc_hd__buf_8 _28853_ (.A(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__a22oi_4 _28854_ (.A1(_05174_),
    .A2(net466),
    .B1(_05142_),
    .B2(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__buf_4 _28855_ (.A(_05235_),
    .X(_06314_));
 sky130_fd_sc_hd__and4_4 _28856_ (.A(_06314_),
    .B(_19934_),
    .C(_06143_),
    .D(_06151_),
    .X(_06315_));
 sky130_fd_sc_hd__nor2_1 _28857_ (.A(_06313_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__o21ai_2 _28858_ (.A1(_05154_),
    .A2(_06308_),
    .B1(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__nor2_1 _28859_ (.A(_05154_),
    .B(_06308_),
    .Y(_06318_));
 sky130_fd_sc_hd__o21ai_2 _28860_ (.A1(_06313_),
    .A2(_06315_),
    .B1(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand2_2 _28861_ (.A(_06317_),
    .B(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__a21o_2 _28862_ (.A1(_06302_),
    .A2(_06306_),
    .B1(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__nand3_4 _28863_ (.A(_06320_),
    .B(_06306_),
    .C(_06302_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2_2 _28864_ (.A(_06175_),
    .B(_06166_),
    .Y(_06323_));
 sky130_fd_sc_hd__a21o_2 _28865_ (.A1(_06321_),
    .A2(_06322_),
    .B1(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__nor2_4 _28866_ (.A(_06157_),
    .B(_06160_),
    .Y(_06325_));
 sky130_fd_sc_hd__nor2_2 _28867_ (.A(_06156_),
    .B(_06325_),
    .Y(_06326_));
 sky130_vsdinv _28868_ (.A(_06326_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand3_4 _28869_ (.A(_06321_),
    .B(_06323_),
    .C(_06322_),
    .Y(_06328_));
 sky130_fd_sc_hd__and3_1 _28870_ (.A(_06324_),
    .B(_06327_),
    .C(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__a21oi_4 _28871_ (.A1(_06324_),
    .A2(_06328_),
    .B1(_06327_),
    .Y(_06330_));
 sky130_fd_sc_hd__o2bb2ai_4 _28872_ (.A1_N(_06282_),
    .A2_N(_06286_),
    .B1(_06329_),
    .B2(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__a21oi_2 _28873_ (.A1(_06321_),
    .A2(_06322_),
    .B1(_06323_),
    .Y(_06332_));
 sky130_fd_sc_hd__o211a_2 _28874_ (.A1(_06162_),
    .A2(_06174_),
    .B1(_06322_),
    .C1(_06321_),
    .X(_06333_));
 sky130_fd_sc_hd__o22ai_4 _28875_ (.A1(_06156_),
    .A2(_06325_),
    .B1(_06332_),
    .B2(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__nand3_4 _28876_ (.A(_06324_),
    .B(_06326_),
    .C(_06328_),
    .Y(_06335_));
 sky130_fd_sc_hd__nand2_2 _28877_ (.A(_06334_),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__nand3_4 _28878_ (.A(_06336_),
    .B(_06282_),
    .C(_06286_),
    .Y(_06337_));
 sky130_vsdinv _28879_ (.A(_06136_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _28880_ (.A(_06132_),
    .B(_06025_),
    .Y(_06339_));
 sky130_fd_sc_hd__o22ai_4 _28881_ (.A1(_06338_),
    .A2(_06339_),
    .B1(_06187_),
    .B2(_06137_),
    .Y(_06340_));
 sky130_fd_sc_hd__a21oi_4 _28882_ (.A1(_06331_),
    .A2(_06337_),
    .B1(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand3_4 _28883_ (.A(_06340_),
    .B(_06337_),
    .C(_06331_),
    .Y(_06342_));
 sky130_fd_sc_hd__a22oi_4 _28884_ (.A1(_06048_),
    .A2(_05183_),
    .B1(_06049_),
    .B2(_05238_),
    .Y(_06343_));
 sky130_fd_sc_hd__buf_6 _28885_ (.A(_06117_),
    .X(_06344_));
 sky130_fd_sc_hd__nand2_2 _28886_ (.A(_06344_),
    .B(_20168_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _28887_ (.A(_06045_),
    .B(_20165_),
    .Y(_06346_));
 sky130_fd_sc_hd__nor2_1 _28888_ (.A(_06345_),
    .B(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__buf_6 _28889_ (.A(_05392_),
    .X(_06348_));
 sky130_fd_sc_hd__nand2_2 _28890_ (.A(_06052_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__o21bai_1 _28891_ (.A1(_06343_),
    .A2(_06347_),
    .B1_N(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand3b_2 _28892_ (.A_N(_06345_),
    .B(_06046_),
    .C(_20166_),
    .Y(_06351_));
 sky130_fd_sc_hd__nand2_1 _28893_ (.A(_06345_),
    .B(_06346_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand3_1 _28894_ (.A(_06351_),
    .B(_06349_),
    .C(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__nand2_2 _28895_ (.A(_06350_),
    .B(_06353_),
    .Y(_06354_));
 sky130_vsdinv _28896_ (.A(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__buf_4 _28897_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06356_));
 sky130_fd_sc_hd__buf_6 _28898_ (.A(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__buf_6 _28899_ (.A(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__buf_8 _28900_ (.A(_19895_),
    .X(_06359_));
 sky130_fd_sc_hd__buf_6 _28901_ (.A(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__a22oi_4 _28902_ (.A1(_06358_),
    .A2(_05415_),
    .B1(_06360_),
    .B2(_05147_),
    .Y(_06361_));
 sky130_fd_sc_hd__nand2_2 _28903_ (.A(_06207_),
    .B(_05297_),
    .Y(_06362_));
 sky130_fd_sc_hd__buf_6 _28904_ (.A(_06356_),
    .X(_06363_));
 sky130_fd_sc_hd__nand2_1 _28905_ (.A(_06363_),
    .B(_04838_),
    .Y(_06364_));
 sky130_fd_sc_hd__nor2_2 _28906_ (.A(_06362_),
    .B(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__clkbuf_4 _28907_ (.A(\pcpi_mul.rs2[12] ),
    .X(_06366_));
 sky130_fd_sc_hd__nand2_2 _28908_ (.A(_06366_),
    .B(_05300_),
    .Y(_06367_));
 sky130_fd_sc_hd__o21bai_2 _28909_ (.A1(_06361_),
    .A2(_06365_),
    .B1_N(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__clkbuf_2 _28910_ (.A(_19893_),
    .X(_06369_));
 sky130_fd_sc_hd__nand3b_4 _28911_ (.A_N(_06362_),
    .B(net444),
    .C(_05415_),
    .Y(_06370_));
 sky130_fd_sc_hd__nand2_2 _28912_ (.A(_06362_),
    .B(_06364_),
    .Y(_06371_));
 sky130_fd_sc_hd__nand3_4 _28913_ (.A(_06370_),
    .B(_06367_),
    .C(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__a21o_2 _28914_ (.A1(_06368_),
    .A2(_06372_),
    .B1(_06211_),
    .X(_06373_));
 sky130_fd_sc_hd__nand3_4 _28915_ (.A(_06368_),
    .B(_06372_),
    .C(_06211_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_2 _28916_ (.A(_06373_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__or2_2 _28917_ (.A(_06355_),
    .B(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__nand2_2 _28918_ (.A(_06375_),
    .B(_06355_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_4 _28919_ (.A(_06376_),
    .B(_06377_),
    .Y(_06378_));
 sky130_vsdinv _28920_ (.A(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_2 _28921_ (.A(_06342_),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__or2_2 _28922_ (.A(_06341_),
    .B(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__nand2_1 _28923_ (.A(_06331_),
    .B(_06337_),
    .Y(_06382_));
 sky130_fd_sc_hd__o21a_1 _28924_ (.A1(_06187_),
    .A2(_06137_),
    .B1(_06188_),
    .X(_06383_));
 sky130_fd_sc_hd__nand2_2 _28925_ (.A(_06382_),
    .B(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_2 _28926_ (.A(_06384_),
    .B(_06342_),
    .Y(_06385_));
 sky130_fd_sc_hd__a21oi_4 _28927_ (.A1(_06385_),
    .A2(_06378_),
    .B1(_06219_),
    .Y(_06386_));
 sky130_fd_sc_hd__nand2_1 _28928_ (.A(_06381_),
    .B(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__a22oi_4 _28929_ (.A1(_06376_),
    .A2(_06377_),
    .B1(_06384_),
    .B2(_06342_),
    .Y(_06388_));
 sky130_fd_sc_hd__nor2_8 _28930_ (.A(_06341_),
    .B(_06380_),
    .Y(_06389_));
 sky130_fd_sc_hd__o22ai_4 _28931_ (.A1(_06216_),
    .A2(_06194_),
    .B1(_06388_),
    .B2(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__and2_2 _28932_ (.A(_06183_),
    .B(_06182_),
    .X(_06391_));
 sky130_fd_sc_hd__nor2_8 _28933_ (.A(_06391_),
    .B(_06193_),
    .Y(_06392_));
 sky130_fd_sc_hd__and2_1 _28934_ (.A(_06193_),
    .B(_06391_),
    .X(_06393_));
 sky130_fd_sc_hd__nor2_4 _28935_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_vsdinv _28936_ (.A(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand3_2 _28937_ (.A(_06387_),
    .B(_06390_),
    .C(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__a21o_1 _28938_ (.A1(_06387_),
    .A2(_06390_),
    .B1(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__nand3b_2 _28939_ (.A_N(_06244_),
    .B(_06396_),
    .C(_06397_),
    .Y(_06398_));
 sky130_vsdinv _28940_ (.A(_06222_),
    .Y(_06399_));
 sky130_fd_sc_hd__nor2_2 _28941_ (.A(_06399_),
    .B(_06039_),
    .Y(_06400_));
 sky130_fd_sc_hd__nand2_2 _28942_ (.A(_06398_),
    .B(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__nand2_1 _28943_ (.A(_06397_),
    .B(_06396_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand2_1 _28944_ (.A(_06402_),
    .B(_06244_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_1 _28945_ (.A(_06398_),
    .B(_06403_),
    .Y(_06404_));
 sky130_vsdinv _28946_ (.A(_06400_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _28947_ (.A(_06229_),
    .B(_06068_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_1 _28948_ (.A(_06406_),
    .B(_06236_),
    .Y(_06407_));
 sky130_fd_sc_hd__a21boi_2 _28949_ (.A1(_06404_),
    .A2(_06405_),
    .B1_N(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _28950_ (.A(_06404_),
    .B(_06405_),
    .Y(_06409_));
 sky130_fd_sc_hd__a21oi_1 _28951_ (.A1(_06409_),
    .A2(_06401_),
    .B1(_06407_),
    .Y(_06410_));
 sky130_fd_sc_hd__a21oi_2 _28952_ (.A1(_06401_),
    .A2(_06408_),
    .B1(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__o22ai_2 _28953_ (.A1(_06230_),
    .A2(_06239_),
    .B1(_06242_),
    .B2(_06243_),
    .Y(_06412_));
 sky130_fd_sc_hd__or2_1 _28954_ (.A(_06411_),
    .B(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__nand2_2 _28955_ (.A(_06412_),
    .B(_06411_),
    .Y(_06414_));
 sky130_fd_sc_hd__and2_1 _28956_ (.A(_06413_),
    .B(_06414_),
    .X(_02633_));
 sky130_fd_sc_hd__nand2_2 _28957_ (.A(_06408_),
    .B(_06401_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand2_2 _28958_ (.A(_06401_),
    .B(_06403_),
    .Y(_06416_));
 sky130_fd_sc_hd__a21oi_4 _28959_ (.A1(_06324_),
    .A2(_06327_),
    .B1(_06333_),
    .Y(_06417_));
 sky130_vsdinv _28960_ (.A(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__and2_2 _28961_ (.A(_06342_),
    .B(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__nor2_8 _28962_ (.A(_06418_),
    .B(_06342_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_2 _28963_ (.A(_05302_),
    .B(_20145_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand2_2 _28964_ (.A(_19924_),
    .B(_05998_),
    .Y(_06422_));
 sky130_fd_sc_hd__nor2_4 _28965_ (.A(_06421_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__and2_1 _28966_ (.A(_06421_),
    .B(_06422_),
    .X(_06424_));
 sky130_fd_sc_hd__nand2_2 _28967_ (.A(_05307_),
    .B(net473),
    .Y(_06425_));
 sky130_vsdinv _28968_ (.A(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__o21ai_2 _28969_ (.A1(_06423_),
    .A2(_06424_),
    .B1(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__or2_2 _28970_ (.A(_06421_),
    .B(_06422_),
    .X(_06428_));
 sky130_fd_sc_hd__nand2_1 _28971_ (.A(_06421_),
    .B(_06422_),
    .Y(_06429_));
 sky130_fd_sc_hd__nand3_2 _28972_ (.A(_06428_),
    .B(_06429_),
    .C(_06425_),
    .Y(_06430_));
 sky130_fd_sc_hd__a2bb2oi_2 _28973_ (.A1_N(_06298_),
    .A2_N(_06290_),
    .B1(_06299_),
    .B2(_06291_),
    .Y(_06431_));
 sky130_fd_sc_hd__nand3_4 _28974_ (.A(_06427_),
    .B(_06430_),
    .C(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__nand2_2 _28975_ (.A(_06426_),
    .B(_06429_),
    .Y(_06433_));
 sky130_fd_sc_hd__o2bb2ai_2 _28976_ (.A1_N(_06291_),
    .A2_N(_06299_),
    .B1(_06288_),
    .B2(_06290_),
    .Y(_06434_));
 sky130_fd_sc_hd__o21ai_2 _28977_ (.A1(_06423_),
    .A2(_06424_),
    .B1(_06425_),
    .Y(_06435_));
 sky130_fd_sc_hd__o211ai_4 _28978_ (.A1(_06423_),
    .A2(_06433_),
    .B1(_06434_),
    .C1(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__buf_6 _28979_ (.A(_06293_),
    .X(_06437_));
 sky130_fd_sc_hd__buf_6 _28980_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06438_));
 sky130_fd_sc_hd__and4_4 _28981_ (.A(_05282_),
    .B(_05477_),
    .C(_06437_),
    .D(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__clkinv_8 _28982_ (.A(_20132_),
    .Y(_06440_));
 sky130_fd_sc_hd__buf_6 _28983_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06441_));
 sky130_fd_sc_hd__buf_6 _28984_ (.A(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__nand2_2 _28985_ (.A(_05282_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__o21a_2 _28986_ (.A1(_05250_),
    .A2(_06440_),
    .B1(_06443_),
    .X(_06444_));
 sky130_vsdinv _28987_ (.A(\pcpi_mul.rs1[12] ),
    .Y(_06445_));
 sky130_fd_sc_hd__clkbuf_4 _28988_ (.A(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__nor2_2 _28989_ (.A(_05153_),
    .B(net465),
    .Y(_06447_));
 sky130_vsdinv _28990_ (.A(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__nor3_4 _28991_ (.A(_06439_),
    .B(_06444_),
    .C(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__o21a_1 _28992_ (.A1(_06439_),
    .A2(_06444_),
    .B1(_06448_),
    .X(_06450_));
 sky130_fd_sc_hd__o2bb2ai_4 _28993_ (.A1_N(_06432_),
    .A2_N(_06436_),
    .B1(_06449_),
    .B2(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__buf_6 _28994_ (.A(_06440_),
    .X(_06452_));
 sky130_fd_sc_hd__o21ai_2 _28995_ (.A1(_05250_),
    .A2(_06452_),
    .B1(_06443_),
    .Y(_06453_));
 sky130_fd_sc_hd__nand3b_1 _28996_ (.A_N(_06439_),
    .B(_06448_),
    .C(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__o21ai_1 _28997_ (.A1(_06439_),
    .A2(_06444_),
    .B1(_06447_),
    .Y(_06455_));
 sky130_fd_sc_hd__nand2_2 _28998_ (.A(_06454_),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand3_4 _28999_ (.A(_06456_),
    .B(_06436_),
    .C(_06432_),
    .Y(_06457_));
 sky130_fd_sc_hd__nand2_4 _29000_ (.A(_06322_),
    .B(_06302_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21o_1 _29001_ (.A1(_06451_),
    .A2(_06457_),
    .B1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__nand3_4 _29002_ (.A(_06458_),
    .B(_06457_),
    .C(_06451_),
    .Y(_06460_));
 sky130_fd_sc_hd__and2_1 _29003_ (.A(_06316_),
    .B(_06318_),
    .X(_06461_));
 sky130_fd_sc_hd__nor2_4 _29004_ (.A(_06315_),
    .B(_06461_),
    .Y(_06462_));
 sky130_vsdinv _29005_ (.A(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__nand3_4 _29006_ (.A(_06459_),
    .B(_06460_),
    .C(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__a21oi_4 _29007_ (.A1(_06451_),
    .A2(_06457_),
    .B1(_06458_),
    .Y(_06465_));
 sky130_vsdinv _29008_ (.A(_06302_),
    .Y(_06466_));
 sky130_fd_sc_hd__a32oi_2 _29009_ (.A1(_06303_),
    .A2(_06304_),
    .A3(_06305_),
    .B1(_06317_),
    .B2(_06319_),
    .Y(_06467_));
 sky130_fd_sc_hd__o211a_1 _29010_ (.A1(_06466_),
    .A2(_06467_),
    .B1(_06457_),
    .C1(_06451_),
    .X(_06468_));
 sky130_fd_sc_hd__o21ai_2 _29011_ (.A1(_06465_),
    .A2(_06468_),
    .B1(_06462_),
    .Y(_06469_));
 sky130_fd_sc_hd__nor2_2 _29012_ (.A(_06272_),
    .B(_06268_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand2_2 _29013_ (.A(_06263_),
    .B(_06245_),
    .Y(_06471_));
 sky130_fd_sc_hd__buf_4 _29014_ (.A(_20154_),
    .X(_06472_));
 sky130_fd_sc_hd__buf_6 _29015_ (.A(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__buf_6 _29016_ (.A(_19914_),
    .X(_06474_));
 sky130_fd_sc_hd__buf_4 _29017_ (.A(\pcpi_mul.rs1[8] ),
    .X(_06475_));
 sky130_fd_sc_hd__buf_6 _29018_ (.A(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__a22oi_4 _29019_ (.A1(_06100_),
    .A2(_06473_),
    .B1(_06474_),
    .B2(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__buf_4 _29020_ (.A(_05501_),
    .X(_06478_));
 sky130_fd_sc_hd__and4_4 _29021_ (.A(_06478_),
    .B(_05499_),
    .C(_05698_),
    .D(_05799_),
    .X(_06479_));
 sky130_fd_sc_hd__buf_6 _29022_ (.A(_05554_),
    .X(_06480_));
 sky130_fd_sc_hd__nand2_2 _29023_ (.A(_19917_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__o21ai_2 _29024_ (.A1(_06477_),
    .A2(_06479_),
    .B1(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__buf_6 _29025_ (.A(_05501_),
    .X(_06483_));
 sky130_fd_sc_hd__nand2_1 _29026_ (.A(_06483_),
    .B(_05573_),
    .Y(_06484_));
 sky130_fd_sc_hd__nand3b_4 _29027_ (.A_N(_06484_),
    .B(_06098_),
    .C(_05832_),
    .Y(_06485_));
 sky130_vsdinv _29028_ (.A(_06481_),
    .Y(_06486_));
 sky130_fd_sc_hd__a22o_2 _29029_ (.A1(_06100_),
    .A2(_06473_),
    .B1(_06474_),
    .B2(_05991_),
    .X(_06487_));
 sky130_fd_sc_hd__nand3_4 _29030_ (.A(_06485_),
    .B(_06486_),
    .C(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__o21ai_2 _29031_ (.A1(_06349_),
    .A2(_06343_),
    .B1(_06351_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand3_4 _29032_ (.A(_06482_),
    .B(_06488_),
    .C(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__o21ai_2 _29033_ (.A1(_06477_),
    .A2(_06479_),
    .B1(_06486_),
    .Y(_06491_));
 sky130_fd_sc_hd__nand3_2 _29034_ (.A(_06485_),
    .B(_06481_),
    .C(_06487_),
    .Y(_06492_));
 sky130_fd_sc_hd__o21ai_1 _29035_ (.A1(_06345_),
    .A2(_06346_),
    .B1(_06349_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_1 _29036_ (.A(_06493_),
    .B(_06352_),
    .Y(_06494_));
 sky130_fd_sc_hd__nand3_4 _29037_ (.A(_06491_),
    .B(_06492_),
    .C(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__nor2_8 _29038_ (.A(_06253_),
    .B(_06251_),
    .Y(_06496_));
 sky130_fd_sc_hd__nor2_4 _29039_ (.A(_06246_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__a21oi_2 _29040_ (.A1(_06490_),
    .A2(_06495_),
    .B1(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__and3_1 _29041_ (.A(_06490_),
    .B(_06495_),
    .C(_06497_),
    .X(_06499_));
 sky130_fd_sc_hd__nand2_1 _29042_ (.A(_06374_),
    .B(_06354_),
    .Y(_06500_));
 sky130_fd_sc_hd__nand2_4 _29043_ (.A(_06500_),
    .B(_06373_),
    .Y(_06501_));
 sky130_fd_sc_hd__o21bai_4 _29044_ (.A1(_06498_),
    .A2(_06499_),
    .B1_N(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__o2bb2ai_4 _29045_ (.A1_N(_06490_),
    .A2_N(_06495_),
    .B1(_06246_),
    .B2(_06496_),
    .Y(_06503_));
 sky130_fd_sc_hd__nand3_4 _29046_ (.A(_06490_),
    .B(_06495_),
    .C(_06497_),
    .Y(_06504_));
 sky130_fd_sc_hd__nand3_4 _29047_ (.A(_06501_),
    .B(_06503_),
    .C(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__a22oi_4 _29048_ (.A1(_06259_),
    .A2(_06471_),
    .B1(_06502_),
    .B2(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand2_4 _29049_ (.A(_06471_),
    .B(_06259_),
    .Y(_06507_));
 sky130_fd_sc_hd__a21oi_4 _29050_ (.A1(_06503_),
    .A2(_06504_),
    .B1(_06501_),
    .Y(_06508_));
 sky130_fd_sc_hd__and3_1 _29051_ (.A(_06482_),
    .B(_06488_),
    .C(_06489_),
    .X(_06509_));
 sky130_fd_sc_hd__nand2_1 _29052_ (.A(_06495_),
    .B(_06497_),
    .Y(_06510_));
 sky130_fd_sc_hd__o211a_2 _29053_ (.A1(_06509_),
    .A2(_06510_),
    .B1(_06503_),
    .C1(_06501_),
    .X(_06511_));
 sky130_fd_sc_hd__nor3_4 _29054_ (.A(_06507_),
    .B(_06508_),
    .C(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__o22ai_4 _29055_ (.A1(_06270_),
    .A2(_06470_),
    .B1(_06506_),
    .B2(_06512_),
    .Y(_06513_));
 sky130_fd_sc_hd__o21ai_4 _29056_ (.A1(_06508_),
    .A2(_06511_),
    .B1(_06507_),
    .Y(_06514_));
 sky130_fd_sc_hd__o21ai_4 _29057_ (.A1(_06280_),
    .A2(_06270_),
    .B1(_06276_),
    .Y(_06515_));
 sky130_fd_sc_hd__nand3b_4 _29058_ (.A_N(_06507_),
    .B(_06502_),
    .C(_06505_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand3_4 _29059_ (.A(_06514_),
    .B(_06515_),
    .C(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__a22oi_4 _29060_ (.A1(_06464_),
    .A2(_06469_),
    .B1(_06513_),
    .B2(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_2 _29061_ (.A(_06514_),
    .B(_06515_),
    .Y(_06519_));
 sky130_fd_sc_hd__o21ai_1 _29062_ (.A1(_06465_),
    .A2(_06468_),
    .B1(_06463_),
    .Y(_06520_));
 sky130_fd_sc_hd__nand3_1 _29063_ (.A(_06459_),
    .B(_06460_),
    .C(_06462_),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_2 _29064_ (.A(_06520_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__o211a_1 _29065_ (.A1(_06512_),
    .A2(_06519_),
    .B1(_06522_),
    .C1(_06513_),
    .X(_06523_));
 sky130_vsdinv _29066_ (.A(_06286_),
    .Y(_06524_));
 sky130_fd_sc_hd__a32oi_4 _29067_ (.A1(_06273_),
    .A2(_06281_),
    .A3(_06275_),
    .B1(_06335_),
    .B2(_06334_),
    .Y(_06525_));
 sky130_fd_sc_hd__nor2_8 _29068_ (.A(_06524_),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__o21ai_4 _29069_ (.A1(_06518_),
    .A2(_06523_),
    .B1(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__clkinv_8 _29070_ (.A(_19889_),
    .Y(_06528_));
 sky130_fd_sc_hd__buf_4 _29071_ (.A(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__nor2_8 _29072_ (.A(_06529_),
    .B(net449),
    .Y(_06530_));
 sky130_fd_sc_hd__buf_8 _29073_ (.A(_06041_),
    .X(_06531_));
 sky130_fd_sc_hd__a22oi_4 _29074_ (.A1(_06531_),
    .A2(_20165_),
    .B1(_06196_),
    .B2(_05481_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand2_1 _29075_ (.A(_06041_),
    .B(_05237_),
    .Y(_06533_));
 sky130_fd_sc_hd__buf_6 _29076_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06534_));
 sky130_fd_sc_hd__nand2_1 _29077_ (.A(_06534_),
    .B(_05388_),
    .Y(_06535_));
 sky130_fd_sc_hd__nor2_1 _29078_ (.A(_06533_),
    .B(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_2 _29079_ (.A(_19909_),
    .B(_06249_),
    .Y(_06537_));
 sky130_fd_sc_hd__o21bai_1 _29080_ (.A1(_06532_),
    .A2(_06536_),
    .B1_N(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__nand3b_2 _29081_ (.A_N(_06533_),
    .B(_06107_),
    .C(_06348_),
    .Y(_06539_));
 sky130_fd_sc_hd__nand2_1 _29082_ (.A(_06533_),
    .B(_06535_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand3_1 _29083_ (.A(_06539_),
    .B(_06540_),
    .C(_06537_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_2 _29084_ (.A(_06538_),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__buf_6 _29085_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_8 _29086_ (.A(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__buf_6 _29087_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06545_));
 sky130_fd_sc_hd__buf_8 _29088_ (.A(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__a22oi_1 _29089_ (.A1(_06544_),
    .A2(_05146_),
    .B1(_06546_),
    .B2(_06197_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand2_4 _29090_ (.A(_06543_),
    .B(_05145_),
    .Y(_06548_));
 sky130_fd_sc_hd__nand2_2 _29091_ (.A(_06545_),
    .B(_05178_),
    .Y(_06549_));
 sky130_fd_sc_hd__nor2_1 _29092_ (.A(_06548_),
    .B(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__buf_6 _29093_ (.A(_20167_),
    .X(_06551_));
 sky130_fd_sc_hd__nand2_2 _29094_ (.A(_06366_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__o21bai_1 _29095_ (.A1(_06547_),
    .A2(_06550_),
    .B1_N(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__nand3b_2 _29096_ (.A_N(_06548_),
    .B(_06208_),
    .C(_05181_),
    .Y(_06554_));
 sky130_fd_sc_hd__nand2_4 _29097_ (.A(_06548_),
    .B(_06549_),
    .Y(_06555_));
 sky130_fd_sc_hd__nand3_2 _29098_ (.A(_06554_),
    .B(_06555_),
    .C(_06552_),
    .Y(_06556_));
 sky130_vsdinv _29099_ (.A(_06367_),
    .Y(_06557_));
 sky130_fd_sc_hd__a21oi_2 _29100_ (.A1(_06557_),
    .A2(_06371_),
    .B1(_06365_),
    .Y(_06558_));
 sky130_fd_sc_hd__a21o_1 _29101_ (.A1(_06553_),
    .A2(_06556_),
    .B1(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__nand3_2 _29102_ (.A(_06553_),
    .B(_06556_),
    .C(_06558_),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_2 _29103_ (.A(_06559_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__xnor2_4 _29104_ (.A(_06542_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__nor2_4 _29105_ (.A(_06530_),
    .B(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__and2_1 _29106_ (.A(_06562_),
    .B(_06530_),
    .X(_06564_));
 sky130_fd_sc_hd__clkbuf_4 _29107_ (.A(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__nor2_4 _29108_ (.A(_06563_),
    .B(_06565_),
    .Y(_06566_));
 sky130_vsdinv _29109_ (.A(_06464_),
    .Y(_06567_));
 sky130_fd_sc_hd__a21oi_2 _29110_ (.A1(_06459_),
    .A2(_06460_),
    .B1(_06463_),
    .Y(_06568_));
 sky130_fd_sc_hd__a21oi_4 _29111_ (.A1(_06514_),
    .A2(_06516_),
    .B1(_06515_),
    .Y(_06569_));
 sky130_fd_sc_hd__a21oi_1 _29112_ (.A1(_06277_),
    .A2(_06278_),
    .B1(_06280_),
    .Y(_06570_));
 sky130_fd_sc_hd__o211a_1 _29113_ (.A1(_06268_),
    .A2(_06570_),
    .B1(_06516_),
    .C1(_06514_),
    .X(_06571_));
 sky130_fd_sc_hd__o22ai_4 _29114_ (.A1(_06567_),
    .A2(_06568_),
    .B1(_06569_),
    .B2(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__nand2_1 _29115_ (.A(_06336_),
    .B(_06282_),
    .Y(_06573_));
 sky130_fd_sc_hd__nand2_2 _29116_ (.A(_06573_),
    .B(_06286_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand3_4 _29117_ (.A(_06513_),
    .B(_06517_),
    .C(_06522_),
    .Y(_06575_));
 sky130_fd_sc_hd__nand3_4 _29118_ (.A(_06572_),
    .B(_06574_),
    .C(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__nand3_4 _29119_ (.A(_06527_),
    .B(_06566_),
    .C(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__a21oi_2 _29120_ (.A1(_06572_),
    .A2(_06575_),
    .B1(_06574_),
    .Y(_06578_));
 sky130_fd_sc_hd__o211a_2 _29121_ (.A1(_06524_),
    .A2(_06525_),
    .B1(_06575_),
    .C1(_06572_),
    .X(_06579_));
 sky130_fd_sc_hd__o22ai_4 _29122_ (.A1(_06565_),
    .A2(_06563_),
    .B1(_06578_),
    .B2(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__a2bb2oi_4 _29123_ (.A1_N(_06385_),
    .A2_N(_06378_),
    .B1(_06577_),
    .B2(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand2_2 _29124_ (.A(_06527_),
    .B(_06566_),
    .Y(_06582_));
 sky130_fd_sc_hd__o211a_2 _29125_ (.A1(_06579_),
    .A2(_06582_),
    .B1(_06389_),
    .C1(_06580_),
    .X(_06583_));
 sky130_fd_sc_hd__o22ai_4 _29126_ (.A1(_06419_),
    .A2(_06420_),
    .B1(_06581_),
    .B2(_06583_),
    .Y(_06584_));
 sky130_fd_sc_hd__a21o_1 _29127_ (.A1(_06580_),
    .A2(_06577_),
    .B1(_06389_),
    .X(_06585_));
 sky130_fd_sc_hd__nand3_4 _29128_ (.A(_06580_),
    .B(_06389_),
    .C(_06577_),
    .Y(_06586_));
 sky130_fd_sc_hd__nor2_8 _29129_ (.A(_06420_),
    .B(_06419_),
    .Y(_06587_));
 sky130_fd_sc_hd__nand3_2 _29130_ (.A(_06585_),
    .B(_06586_),
    .C(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__a22oi_4 _29131_ (.A1(_06381_),
    .A2(_06386_),
    .B1(_06390_),
    .B2(_06394_),
    .Y(_06589_));
 sky130_fd_sc_hd__nand3_4 _29132_ (.A(_06584_),
    .B(_06588_),
    .C(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__nor3_4 _29133_ (.A(_06587_),
    .B(_06581_),
    .C(_06583_),
    .Y(_06591_));
 sky130_fd_sc_hd__a22o_1 _29134_ (.A1(_06381_),
    .A2(_06386_),
    .B1(_06390_),
    .B2(_06394_),
    .X(_06592_));
 sky130_fd_sc_hd__o21ai_1 _29135_ (.A1(_06581_),
    .A2(_06583_),
    .B1(_06587_),
    .Y(_06593_));
 sky130_fd_sc_hd__nand2_1 _29136_ (.A(_06592_),
    .B(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__or2_1 _29137_ (.A(_06591_),
    .B(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__a21o_1 _29138_ (.A1(_06595_),
    .A2(_06590_),
    .B1(_06392_),
    .X(_06596_));
 sky130_fd_sc_hd__a21boi_4 _29139_ (.A1(_06392_),
    .A2(_06590_),
    .B1_N(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__nor2_1 _29140_ (.A(_06416_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand2_1 _29141_ (.A(_06597_),
    .B(_06416_),
    .Y(_06599_));
 sky130_fd_sc_hd__nand3_4 _29142_ (.A(_06414_),
    .B(_06415_),
    .C(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__o21a_2 _29143_ (.A1(_06597_),
    .A2(_06416_),
    .B1(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__a31oi_1 _29144_ (.A1(_06415_),
    .A2(_06414_),
    .A3(_06598_),
    .B1(_06601_),
    .Y(_02634_));
 sky130_fd_sc_hd__o21a_2 _29145_ (.A1(_06462_),
    .A2(_06465_),
    .B1(_06460_),
    .X(_06602_));
 sky130_fd_sc_hd__nor2_4 _29146_ (.A(_06602_),
    .B(_06576_),
    .Y(_06603_));
 sky130_fd_sc_hd__and2_1 _29147_ (.A(_06576_),
    .B(_06602_),
    .X(_06604_));
 sky130_fd_sc_hd__nor2_2 _29148_ (.A(_06603_),
    .B(_06604_),
    .Y(_06605_));
 sky130_fd_sc_hd__buf_4 _29149_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06606_));
 sky130_fd_sc_hd__buf_8 _29150_ (.A(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__a22oi_4 _29151_ (.A1(_06363_),
    .A2(_05143_),
    .B1(_06607_),
    .B2(_05451_),
    .Y(_06608_));
 sky130_fd_sc_hd__nand2_4 _29152_ (.A(_19892_),
    .B(_05299_),
    .Y(_06609_));
 sky130_fd_sc_hd__nand2_4 _29153_ (.A(_06545_),
    .B(_05602_),
    .Y(_06610_));
 sky130_fd_sc_hd__nor2_8 _29154_ (.A(_06609_),
    .B(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__nand2_4 _29155_ (.A(_19898_),
    .B(_05460_),
    .Y(_06612_));
 sky130_fd_sc_hd__o21bai_2 _29156_ (.A1(_06608_),
    .A2(_06611_),
    .B1_N(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__buf_6 _29157_ (.A(_05602_),
    .X(_06614_));
 sky130_fd_sc_hd__nand3b_4 _29158_ (.A_N(_06609_),
    .B(_06546_),
    .C(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_2 _29159_ (.A(_06609_),
    .B(_06610_),
    .Y(_06616_));
 sky130_fd_sc_hd__nand3_4 _29160_ (.A(_06615_),
    .B(_06612_),
    .C(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__o21ai_4 _29161_ (.A1(_06548_),
    .A2(_06549_),
    .B1(_06552_),
    .Y(_06618_));
 sky130_fd_sc_hd__nand2_2 _29162_ (.A(_06618_),
    .B(_06555_),
    .Y(_06619_));
 sky130_fd_sc_hd__a21o_1 _29163_ (.A1(_06613_),
    .A2(_06617_),
    .B1(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__nand3_4 _29164_ (.A(_06613_),
    .B(_06617_),
    .C(_06619_),
    .Y(_06621_));
 sky130_fd_sc_hd__buf_4 _29165_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06622_));
 sky130_fd_sc_hd__nand2_8 _29166_ (.A(_06622_),
    .B(_05656_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_8 _29167_ (.A(_05664_),
    .B(_05285_),
    .Y(_06624_));
 sky130_fd_sc_hd__nor2_2 _29168_ (.A(_06623_),
    .B(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__nand2_4 _29169_ (.A(_19908_),
    .B(_06472_),
    .Y(_06626_));
 sky130_fd_sc_hd__buf_4 _29170_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06627_));
 sky130_fd_sc_hd__a22o_2 _29171_ (.A1(_06627_),
    .A2(_05218_),
    .B1(_19905_),
    .B2(_05389_),
    .X(_06628_));
 sky130_fd_sc_hd__nand3b_4 _29172_ (.A_N(_06625_),
    .B(_06626_),
    .C(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__buf_8 _29173_ (.A(_06622_),
    .X(_06630_));
 sky130_fd_sc_hd__buf_6 _29174_ (.A(_05656_),
    .X(_06631_));
 sky130_fd_sc_hd__a22oi_4 _29175_ (.A1(_06630_),
    .A2(_05388_),
    .B1(_06631_),
    .B2(_05665_),
    .Y(_06632_));
 sky130_vsdinv _29176_ (.A(_06626_),
    .Y(_06633_));
 sky130_fd_sc_hd__o21ai_2 _29177_ (.A1(_06632_),
    .A2(_06625_),
    .B1(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__nand2_2 _29178_ (.A(_06629_),
    .B(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__buf_4 _29179_ (.A(\pcpi_mul.rs2[16] ),
    .X(_06636_));
 sky130_fd_sc_hd__buf_6 _29180_ (.A(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__buf_6 _29181_ (.A(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__nand2_2 _29182_ (.A(_06638_),
    .B(_05415_),
    .Y(_06639_));
 sky130_fd_sc_hd__buf_6 _29183_ (.A(_19889_),
    .X(_06640_));
 sky130_fd_sc_hd__buf_8 _29184_ (.A(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__nand2_2 _29185_ (.A(_06641_),
    .B(_05147_),
    .Y(_06642_));
 sky130_fd_sc_hd__nor2_2 _29186_ (.A(_06639_),
    .B(_06642_),
    .Y(_06643_));
 sky130_vsdinv _29187_ (.A(_06643_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_1 _29188_ (.A(_06639_),
    .B(_06642_),
    .Y(_06645_));
 sky130_fd_sc_hd__nand2_1 _29189_ (.A(_06644_),
    .B(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__a31o_1 _29190_ (.A1(_06620_),
    .A2(_06621_),
    .A3(_06635_),
    .B1(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__nand2_1 _29191_ (.A(_06620_),
    .B(_06621_),
    .Y(_06648_));
 sky130_vsdinv _29192_ (.A(_06635_),
    .Y(_06649_));
 sky130_fd_sc_hd__nand2_1 _29193_ (.A(_06648_),
    .B(_06649_),
    .Y(_06650_));
 sky130_vsdinv _29194_ (.A(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__or2_4 _29195_ (.A(_06647_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__a21o_1 _29196_ (.A1(_06634_),
    .A2(_06629_),
    .B1(_06648_),
    .X(_06653_));
 sky130_fd_sc_hd__a22o_2 _29197_ (.A1(_06645_),
    .A2(_06644_),
    .B1(_06653_),
    .B2(_06650_),
    .X(_06654_));
 sky130_fd_sc_hd__nand3_4 _29198_ (.A(_06565_),
    .B(_06652_),
    .C(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__a21o_1 _29199_ (.A1(_06652_),
    .A2(_06654_),
    .B1(_06565_),
    .X(_06656_));
 sky130_fd_sc_hd__clkbuf_8 _29200_ (.A(_05724_),
    .X(_06657_));
 sky130_fd_sc_hd__a22oi_4 _29201_ (.A1(_06095_),
    .A2(_05831_),
    .B1(_06657_),
    .B2(_05699_),
    .Y(_06658_));
 sky130_fd_sc_hd__buf_6 _29202_ (.A(\pcpi_mul.rs2[8] ),
    .X(_06659_));
 sky130_fd_sc_hd__nand3_4 _29203_ (.A(_06659_),
    .B(_06110_),
    .C(_06475_),
    .Y(_06660_));
 sky130_fd_sc_hd__nor2_8 _29204_ (.A(_06003_),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_2 _29205_ (.A(_05601_),
    .B(_20145_),
    .Y(_06662_));
 sky130_fd_sc_hd__o21ai_2 _29206_ (.A1(_06658_),
    .A2(_06661_),
    .B1(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__o21ai_2 _29207_ (.A1(_06537_),
    .A2(_06532_),
    .B1(_06539_),
    .Y(_06664_));
 sky130_vsdinv _29208_ (.A(_06662_),
    .Y(_06665_));
 sky130_fd_sc_hd__a22o_1 _29209_ (.A1(_06483_),
    .A2(_05463_),
    .B1(_19915_),
    .B2(_20149_),
    .X(_06666_));
 sky130_fd_sc_hd__o211ai_2 _29210_ (.A1(_06004_),
    .A2(_06660_),
    .B1(_06665_),
    .C1(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand3_4 _29211_ (.A(_06663_),
    .B(_06664_),
    .C(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__o21ai_2 _29212_ (.A1(_06658_),
    .A2(_06661_),
    .B1(_06665_),
    .Y(_06669_));
 sky130_fd_sc_hd__o21ai_1 _29213_ (.A1(_06533_),
    .A2(_06535_),
    .B1(_06537_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand2_1 _29214_ (.A(_06670_),
    .B(_06540_),
    .Y(_06671_));
 sky130_fd_sc_hd__buf_8 _29215_ (.A(_06003_),
    .X(_06672_));
 sky130_fd_sc_hd__o211ai_2 _29216_ (.A1(_06672_),
    .A2(_06660_),
    .B1(_06662_),
    .C1(_06666_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand3_4 _29217_ (.A(_06669_),
    .B(_06671_),
    .C(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__nor2_8 _29218_ (.A(_06486_),
    .B(_06479_),
    .Y(_06675_));
 sky130_fd_sc_hd__o2bb2ai_4 _29219_ (.A1_N(_06668_),
    .A2_N(_06674_),
    .B1(_06477_),
    .B2(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__nor2_4 _29220_ (.A(_06477_),
    .B(_06675_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand3_4 _29221_ (.A(_06668_),
    .B(_06674_),
    .C(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__nand2_1 _29222_ (.A(_06560_),
    .B(_06542_),
    .Y(_06679_));
 sky130_fd_sc_hd__nand2_4 _29223_ (.A(_06679_),
    .B(_06559_),
    .Y(_06680_));
 sky130_fd_sc_hd__a21oi_4 _29224_ (.A1(_06676_),
    .A2(_06678_),
    .B1(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__nand2_1 _29225_ (.A(_06674_),
    .B(_06677_),
    .Y(_06682_));
 sky130_vsdinv _29226_ (.A(_06668_),
    .Y(_06683_));
 sky130_fd_sc_hd__o211a_1 _29227_ (.A1(_06682_),
    .A2(_06683_),
    .B1(_06676_),
    .C1(_06680_),
    .X(_06684_));
 sky130_fd_sc_hd__and2_2 _29228_ (.A(_06510_),
    .B(_06490_),
    .X(_06685_));
 sky130_fd_sc_hd__o21ai_4 _29229_ (.A1(_06681_),
    .A2(_06684_),
    .B1(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__a21o_1 _29230_ (.A1(_06676_),
    .A2(_06678_),
    .B1(_06680_),
    .X(_06687_));
 sky130_fd_sc_hd__nand3_4 _29231_ (.A(_06680_),
    .B(_06676_),
    .C(_06678_),
    .Y(_06688_));
 sky130_fd_sc_hd__nand3b_4 _29232_ (.A_N(_06685_),
    .B(_06687_),
    .C(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__o21ai_4 _29233_ (.A1(_06507_),
    .A2(_06508_),
    .B1(_06505_),
    .Y(_06690_));
 sky130_fd_sc_hd__a21oi_4 _29234_ (.A1(_06686_),
    .A2(_06689_),
    .B1(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__nor2_1 _29235_ (.A(_06507_),
    .B(_06508_),
    .Y(_06692_));
 sky130_fd_sc_hd__o211a_2 _29236_ (.A1(_06511_),
    .A2(_06692_),
    .B1(_06689_),
    .C1(_06686_),
    .X(_06693_));
 sky130_fd_sc_hd__nand2_2 _29237_ (.A(_06428_),
    .B(_06433_),
    .Y(_06694_));
 sky130_fd_sc_hd__buf_6 _29238_ (.A(_06152_),
    .X(_06695_));
 sky130_fd_sc_hd__buf_6 _29239_ (.A(_20137_),
    .X(_06696_));
 sky130_fd_sc_hd__a22oi_4 _29240_ (.A1(_05311_),
    .A2(_06695_),
    .B1(_05312_),
    .B2(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__nand2_4 _29241_ (.A(_19919_),
    .B(_05998_),
    .Y(_06698_));
 sky130_fd_sc_hd__nand2_4 _29242_ (.A(_19924_),
    .B(_05985_),
    .Y(_06699_));
 sky130_fd_sc_hd__nor2_8 _29243_ (.A(_06698_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__buf_6 _29244_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06701_));
 sky130_fd_sc_hd__nand2_2 _29245_ (.A(_05307_),
    .B(_06701_),
    .Y(_06702_));
 sky130_vsdinv _29246_ (.A(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__o21ai_2 _29247_ (.A1(_06697_),
    .A2(_06700_),
    .B1(_06703_),
    .Y(_06704_));
 sky130_vsdinv _29248_ (.A(_06700_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_2 _29249_ (.A(_06698_),
    .B(_06699_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand3_2 _29250_ (.A(_06705_),
    .B(_06702_),
    .C(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__nand3b_4 _29251_ (.A_N(_06694_),
    .B(_06704_),
    .C(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand3_4 _29252_ (.A(_06705_),
    .B(_06703_),
    .C(_06706_),
    .Y(_06709_));
 sky130_fd_sc_hd__o21ai_2 _29253_ (.A1(_06697_),
    .A2(_06700_),
    .B1(_06702_),
    .Y(_06710_));
 sky130_fd_sc_hd__nand3_4 _29254_ (.A(_06709_),
    .B(_06694_),
    .C(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_1 _29255_ (.A(_06708_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__buf_4 _29256_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06713_));
 sky130_fd_sc_hd__buf_6 _29257_ (.A(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__buf_6 _29258_ (.A(_06293_),
    .X(_06715_));
 sky130_fd_sc_hd__nand2_2 _29259_ (.A(_05387_),
    .B(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__a21o_2 _29260_ (.A1(_19934_),
    .A2(_06714_),
    .B1(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__buf_6 _29261_ (.A(_20132_),
    .X(_06718_));
 sky130_fd_sc_hd__buf_4 _29262_ (.A(_20128_),
    .X(_06719_));
 sky130_fd_sc_hd__nand2_2 _29263_ (.A(_05570_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__a21o_1 _29264_ (.A1(_05240_),
    .A2(_06718_),
    .B1(_06720_),
    .X(_06721_));
 sky130_fd_sc_hd__clkinv_8 _29265_ (.A(_06441_),
    .Y(_06722_));
 sky130_fd_sc_hd__nor2_1 _29266_ (.A(_05153_),
    .B(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21bo_2 _29267_ (.A1(_06717_),
    .A2(_06721_),
    .B1_N(_06723_),
    .X(_06724_));
 sky130_vsdinv _29268_ (.A(_06723_),
    .Y(_06725_));
 sky130_fd_sc_hd__nand3_4 _29269_ (.A(_06725_),
    .B(_06717_),
    .C(_06721_),
    .Y(_06726_));
 sky130_fd_sc_hd__and2_1 _29270_ (.A(_06724_),
    .B(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__nand2_1 _29271_ (.A(_06712_),
    .B(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__a21boi_2 _29272_ (.A1(_06456_),
    .A2(_06432_),
    .B1_N(_06436_),
    .Y(_06729_));
 sky130_fd_sc_hd__nand2_2 _29273_ (.A(_06724_),
    .B(_06726_),
    .Y(_06730_));
 sky130_fd_sc_hd__nand3_2 _29274_ (.A(_06708_),
    .B(_06730_),
    .C(_06711_),
    .Y(_06731_));
 sky130_fd_sc_hd__nand3_4 _29275_ (.A(_06728_),
    .B(_06729_),
    .C(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__nand2_2 _29276_ (.A(_06712_),
    .B(_06730_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_2 _29277_ (.A(_06457_),
    .B(_06436_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand3_4 _29278_ (.A(_06727_),
    .B(_06708_),
    .C(_06711_),
    .Y(_06735_));
 sky130_fd_sc_hd__nor2_8 _29279_ (.A(_06439_),
    .B(_06449_),
    .Y(_06736_));
 sky130_fd_sc_hd__a31oi_4 _29280_ (.A1(_06733_),
    .A2(_06734_),
    .A3(_06735_),
    .B1(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand3_4 _29281_ (.A(_06733_),
    .B(_06734_),
    .C(_06735_),
    .Y(_06738_));
 sky130_fd_sc_hd__a21boi_4 _29282_ (.A1(_06738_),
    .A2(_06732_),
    .B1_N(_06736_),
    .Y(_06739_));
 sky130_fd_sc_hd__a21oi_4 _29283_ (.A1(_06732_),
    .A2(_06737_),
    .B1(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__o21ai_2 _29284_ (.A1(_06691_),
    .A2(_06693_),
    .B1(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__a21oi_2 _29285_ (.A1(_06513_),
    .A2(_06522_),
    .B1(_06571_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _29286_ (.A(_06738_),
    .B(_06732_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor2_4 _29287_ (.A(_06736_),
    .B(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__nand3_4 _29288_ (.A(_06686_),
    .B(_06690_),
    .C(_06689_),
    .Y(_06745_));
 sky130_fd_sc_hd__a21o_1 _29289_ (.A1(_06686_),
    .A2(_06689_),
    .B1(_06690_),
    .X(_06746_));
 sky130_fd_sc_hd__o211ai_4 _29290_ (.A1(_06744_),
    .A2(_06739_),
    .B1(_06745_),
    .C1(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__nand3_4 _29291_ (.A(_06741_),
    .B(_06742_),
    .C(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__o22ai_4 _29292_ (.A1(_06744_),
    .A2(_06739_),
    .B1(_06691_),
    .B2(_06693_),
    .Y(_06749_));
 sky130_fd_sc_hd__nand2_1 _29293_ (.A(_06469_),
    .B(_06464_),
    .Y(_06750_));
 sky130_fd_sc_hd__o22ai_4 _29294_ (.A1(_06512_),
    .A2(_06519_),
    .B1(_06750_),
    .B2(_06569_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand3_4 _29295_ (.A(_06746_),
    .B(_06740_),
    .C(_06745_),
    .Y(_06752_));
 sky130_fd_sc_hd__nand3_4 _29296_ (.A(_06749_),
    .B(_06751_),
    .C(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__a22oi_4 _29297_ (.A1(_06655_),
    .A2(_06656_),
    .B1(_06748_),
    .B2(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__nand2_1 _29298_ (.A(_06652_),
    .B(_06654_),
    .Y(_06755_));
 sky130_fd_sc_hd__and2_1 _29299_ (.A(_06755_),
    .B(_06565_),
    .X(_06756_));
 sky130_fd_sc_hd__nor2_1 _29300_ (.A(_06565_),
    .B(_06755_),
    .Y(_06757_));
 sky130_fd_sc_hd__o211a_4 _29301_ (.A1(_06756_),
    .A2(_06757_),
    .B1(_06753_),
    .C1(_06748_),
    .X(_06758_));
 sky130_fd_sc_hd__o22ai_4 _29302_ (.A1(_06579_),
    .A2(_06582_),
    .B1(_06754_),
    .B2(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_2 _29303_ (.A(_06572_),
    .B(_06575_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_2 _29304_ (.A(_06656_),
    .B(_06655_),
    .Y(_06761_));
 sky130_fd_sc_hd__clkbuf_4 _29305_ (.A(_06753_),
    .X(_06762_));
 sky130_fd_sc_hd__nand3b_2 _29306_ (.A_N(_06761_),
    .B(_06748_),
    .C(_06762_),
    .Y(_06763_));
 sky130_fd_sc_hd__a21boi_2 _29307_ (.A1(_06760_),
    .A2(_06526_),
    .B1_N(_06566_),
    .Y(_06764_));
 sky130_fd_sc_hd__and4_1 _29308_ (.A(_06652_),
    .B(_06530_),
    .C(_06654_),
    .D(_06562_),
    .X(_06765_));
 sky130_vsdinv _29309_ (.A(_06656_),
    .Y(_06766_));
 sky130_fd_sc_hd__o2bb2ai_1 _29310_ (.A1_N(_06762_),
    .A2_N(_06748_),
    .B1(_06765_),
    .B2(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__o2111ai_4 _29311_ (.A1(_06526_),
    .A2(_06760_),
    .B1(_06763_),
    .C1(_06764_),
    .D1(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand3b_2 _29312_ (.A_N(_06605_),
    .B(_06759_),
    .C(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__nor2_1 _29313_ (.A(_06602_),
    .B(_06579_),
    .Y(_06770_));
 sky130_fd_sc_hd__and2_1 _29314_ (.A(_06579_),
    .B(_06602_),
    .X(_06771_));
 sky130_fd_sc_hd__o2bb2ai_1 _29315_ (.A1_N(_06768_),
    .A2_N(_06759_),
    .B1(_06770_),
    .B2(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__o2111ai_4 _29316_ (.A1(_06581_),
    .A2(_06587_),
    .B1(_06586_),
    .C1(_06769_),
    .D1(_06772_),
    .Y(_06773_));
 sky130_vsdinv _29317_ (.A(_06577_),
    .Y(_06774_));
 sky130_fd_sc_hd__nand2_1 _29318_ (.A(_06580_),
    .B(_06389_),
    .Y(_06775_));
 sky130_fd_sc_hd__o22ai_4 _29319_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06587_),
    .B2(_06581_),
    .Y(_06776_));
 sky130_fd_sc_hd__o2bb2ai_2 _29320_ (.A1_N(_06768_),
    .A2_N(_06759_),
    .B1(_06603_),
    .B2(_06604_),
    .Y(_06777_));
 sky130_fd_sc_hd__nand3_2 _29321_ (.A(_06759_),
    .B(_06768_),
    .C(_06605_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand3_4 _29322_ (.A(_06776_),
    .B(_06777_),
    .C(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__nor2_4 _29323_ (.A(_06417_),
    .B(_06342_),
    .Y(_06780_));
 sky130_fd_sc_hd__a21oi_1 _29324_ (.A1(_06773_),
    .A2(_06779_),
    .B1(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__and3_1 _29325_ (.A(_06773_),
    .B(_06779_),
    .C(_06780_),
    .X(_06782_));
 sky130_fd_sc_hd__o2bb2ai_2 _29326_ (.A1_N(_06392_),
    .A2_N(_06590_),
    .B1(_06591_),
    .B2(_06594_),
    .Y(_06783_));
 sky130_fd_sc_hd__o21bai_1 _29327_ (.A1(_06781_),
    .A2(_06782_),
    .B1_N(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__a21o_1 _29328_ (.A1(_06773_),
    .A2(_06779_),
    .B1(_06780_),
    .X(_06785_));
 sky130_fd_sc_hd__nand3_4 _29329_ (.A(_06773_),
    .B(_06779_),
    .C(_06780_),
    .Y(_06786_));
 sky130_fd_sc_hd__nand3_4 _29330_ (.A(_06785_),
    .B(_06783_),
    .C(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__nand2_1 _29331_ (.A(_06784_),
    .B(_06787_),
    .Y(_06788_));
 sky130_vsdinv _29332_ (.A(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__nor2_1 _29333_ (.A(_06789_),
    .B(_06601_),
    .Y(_06790_));
 sky130_fd_sc_hd__nand2_1 _29334_ (.A(_06601_),
    .B(_06789_),
    .Y(_06791_));
 sky130_vsdinv _29335_ (.A(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__nor2_1 _29336_ (.A(_06790_),
    .B(_06792_),
    .Y(_02635_));
 sky130_fd_sc_hd__a21bo_2 _29337_ (.A1(_06736_),
    .A2(_06738_),
    .B1_N(_06732_),
    .X(_06793_));
 sky130_fd_sc_hd__nor2_8 _29338_ (.A(_06793_),
    .B(_06762_),
    .Y(_06794_));
 sky130_fd_sc_hd__and2_2 _29339_ (.A(_06762_),
    .B(_06793_),
    .X(_06795_));
 sky130_fd_sc_hd__nor2_8 _29340_ (.A(_06716_),
    .B(_06720_),
    .Y(_06796_));
 sky130_vsdinv _29341_ (.A(_06724_),
    .Y(_06797_));
 sky130_fd_sc_hd__a21oi_2 _29342_ (.A1(_06709_),
    .A2(_06710_),
    .B1(_06694_),
    .Y(_06798_));
 sky130_fd_sc_hd__o21ai_2 _29343_ (.A1(_06730_),
    .A2(_06798_),
    .B1(_06711_),
    .Y(_06799_));
 sky130_fd_sc_hd__nand2_4 _29344_ (.A(_19919_),
    .B(_05985_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_4 _29345_ (.A(_05366_),
    .B(_06441_),
    .Y(_06801_));
 sky130_fd_sc_hd__or2_2 _29346_ (.A(_06800_),
    .B(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__nand2_2 _29347_ (.A(_06800_),
    .B(_06801_),
    .Y(_06803_));
 sky130_fd_sc_hd__nand2_4 _29348_ (.A(_19936_),
    .B(_20122_),
    .Y(_06804_));
 sky130_fd_sc_hd__nand3_2 _29349_ (.A(_06802_),
    .B(_06803_),
    .C(_06804_),
    .Y(_06805_));
 sky130_fd_sc_hd__a21oi_2 _29350_ (.A1(_06703_),
    .A2(_06706_),
    .B1(_06700_),
    .Y(_06806_));
 sky130_fd_sc_hd__a22oi_4 _29351_ (.A1(_05228_),
    .A2(_06696_),
    .B1(_05367_),
    .B2(_06438_),
    .Y(_06807_));
 sky130_fd_sc_hd__nor2_8 _29352_ (.A(_06800_),
    .B(_06801_),
    .Y(_06808_));
 sky130_vsdinv _29353_ (.A(_06804_),
    .Y(_06809_));
 sky130_fd_sc_hd__o21ai_2 _29354_ (.A1(_06807_),
    .A2(_06808_),
    .B1(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand3_4 _29355_ (.A(_06805_),
    .B(_06806_),
    .C(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__nand2_1 _29356_ (.A(_05241_),
    .B(_20125_),
    .Y(_06812_));
 sky130_fd_sc_hd__buf_6 _29357_ (.A(_20128_),
    .X(_06813_));
 sky130_fd_sc_hd__nand3_2 _29358_ (.A(_06812_),
    .B(_05173_),
    .C(_06813_),
    .Y(_06814_));
 sky130_fd_sc_hd__nand2_2 _29359_ (.A(_05235_),
    .B(_06713_),
    .Y(_06815_));
 sky130_fd_sc_hd__buf_6 _29360_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06816_));
 sky130_fd_sc_hd__nand3_4 _29361_ (.A(_06815_),
    .B(_05570_),
    .C(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__nand2_1 _29362_ (.A(_19927_),
    .B(_06437_),
    .Y(_06818_));
 sky130_fd_sc_hd__a21oi_4 _29363_ (.A1(_06814_),
    .A2(_06817_),
    .B1(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__and3_2 _29364_ (.A(_06814_),
    .B(_06817_),
    .C(_06818_),
    .X(_06820_));
 sky130_fd_sc_hd__nor2_4 _29365_ (.A(_06819_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__nand2_2 _29366_ (.A(_06809_),
    .B(_06803_),
    .Y(_06822_));
 sky130_fd_sc_hd__nor2_2 _29367_ (.A(_06702_),
    .B(_06697_),
    .Y(_06823_));
 sky130_fd_sc_hd__o21ai_2 _29368_ (.A1(_06807_),
    .A2(_06808_),
    .B1(_06804_),
    .Y(_06824_));
 sky130_fd_sc_hd__o221ai_4 _29369_ (.A1(_06808_),
    .A2(_06822_),
    .B1(_06700_),
    .B2(_06823_),
    .C1(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__nand3_2 _29370_ (.A(_06811_),
    .B(_06821_),
    .C(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__a21o_1 _29371_ (.A1(_06811_),
    .A2(_06825_),
    .B1(_06821_),
    .X(_06827_));
 sky130_fd_sc_hd__nand3_4 _29372_ (.A(_06799_),
    .B(_06826_),
    .C(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__a21oi_2 _29373_ (.A1(_06811_),
    .A2(_06825_),
    .B1(_06821_),
    .Y(_06829_));
 sky130_fd_sc_hd__and3_1 _29374_ (.A(_06811_),
    .B(_06821_),
    .C(_06825_),
    .X(_06830_));
 sky130_fd_sc_hd__o21a_1 _29375_ (.A1(_06730_),
    .A2(_06798_),
    .B1(_06711_),
    .X(_06831_));
 sky130_fd_sc_hd__o21ai_4 _29376_ (.A1(_06829_),
    .A2(_06830_),
    .B1(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__o211a_4 _29377_ (.A1(_06796_),
    .A2(_06797_),
    .B1(_06828_),
    .C1(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__nor2_1 _29378_ (.A(_06796_),
    .B(_06797_),
    .Y(_06834_));
 sky130_vsdinv _29379_ (.A(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__a21oi_4 _29380_ (.A1(_06832_),
    .A2(_06828_),
    .B1(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_1 _29381_ (.A(_06688_),
    .B(_06685_),
    .Y(_06837_));
 sky130_vsdinv _29382_ (.A(_06674_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_2 _29383_ (.A(_06677_),
    .B(_06683_),
    .Y(_06839_));
 sky130_fd_sc_hd__clkbuf_8 _29384_ (.A(_05412_),
    .X(_06840_));
 sky130_fd_sc_hd__buf_6 _29385_ (.A(_20144_),
    .X(_06841_));
 sky130_fd_sc_hd__a22oi_4 _29386_ (.A1(_05511_),
    .A2(_06480_),
    .B1(_06840_),
    .B2(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__nand3_4 _29387_ (.A(_05722_),
    .B(_05724_),
    .C(_20148_),
    .Y(_06843_));
 sky130_fd_sc_hd__nor2_4 _29388_ (.A(_06287_),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__nand2_2 _29389_ (.A(\pcpi_mul.rs2[6] ),
    .B(_05998_),
    .Y(_06845_));
 sky130_fd_sc_hd__o21ai_2 _29390_ (.A1(_06842_),
    .A2(_06844_),
    .B1(_06845_),
    .Y(_06846_));
 sky130_vsdinv _29391_ (.A(_06845_),
    .Y(_06847_));
 sky130_fd_sc_hd__a22o_1 _29392_ (.A1(_05511_),
    .A2(_06480_),
    .B1(_06840_),
    .B2(_06841_),
    .X(_06848_));
 sky130_fd_sc_hd__o211ai_2 _29393_ (.A1(net445),
    .A2(_06843_),
    .B1(_06847_),
    .C1(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__o22ai_4 _29394_ (.A1(_06623_),
    .A2(_06624_),
    .B1(_06626_),
    .B2(_06632_),
    .Y(_06850_));
 sky130_fd_sc_hd__nand3_4 _29395_ (.A(_06846_),
    .B(_06849_),
    .C(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__o21ai_2 _29396_ (.A1(_06842_),
    .A2(_06844_),
    .B1(_06847_),
    .Y(_06852_));
 sky130_fd_sc_hd__a21oi_2 _29397_ (.A1(_06628_),
    .A2(_06633_),
    .B1(_06625_),
    .Y(_06853_));
 sky130_fd_sc_hd__o211ai_4 _29398_ (.A1(net445),
    .A2(_06843_),
    .B1(_06845_),
    .C1(_06848_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand3_4 _29399_ (.A(_06852_),
    .B(_06853_),
    .C(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__nor2_8 _29400_ (.A(_06665_),
    .B(_06661_),
    .Y(_06856_));
 sky130_fd_sc_hd__o2bb2ai_4 _29401_ (.A1_N(_06851_),
    .A2_N(_06855_),
    .B1(_06658_),
    .B2(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2_4 _29402_ (.A(_06658_),
    .B(_06856_),
    .Y(_06858_));
 sky130_fd_sc_hd__nand3_4 _29403_ (.A(_06855_),
    .B(_06851_),
    .C(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__o21a_1 _29404_ (.A1(_06608_),
    .A2(_06611_),
    .B1(_06612_),
    .X(_06860_));
 sky130_fd_sc_hd__o311ai_4 _29405_ (.A1(_06612_),
    .A2(_06608_),
    .A3(_06611_),
    .B1(_06555_),
    .C1(_06618_),
    .Y(_06861_));
 sky130_fd_sc_hd__o2bb2ai_4 _29406_ (.A1_N(_06621_),
    .A2_N(_06635_),
    .B1(_06860_),
    .B2(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21oi_4 _29407_ (.A1(_06857_),
    .A2(_06859_),
    .B1(_06862_),
    .Y(_06863_));
 sky130_vsdinv _29408_ (.A(_06851_),
    .Y(_06864_));
 sky130_fd_sc_hd__nand2_1 _29409_ (.A(_06855_),
    .B(_06858_),
    .Y(_06865_));
 sky130_fd_sc_hd__o211a_1 _29410_ (.A1(_06864_),
    .A2(_06865_),
    .B1(_06862_),
    .C1(_06857_),
    .X(_06866_));
 sky130_fd_sc_hd__o22ai_4 _29411_ (.A1(_06838_),
    .A2(_06839_),
    .B1(_06863_),
    .B2(_06866_),
    .Y(_06867_));
 sky130_vsdinv _29412_ (.A(_06678_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand3_4 _29413_ (.A(_06857_),
    .B(_06862_),
    .C(_06859_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand2_1 _29414_ (.A(_06857_),
    .B(_06859_),
    .Y(_06870_));
 sky130_fd_sc_hd__o2bb2a_1 _29415_ (.A1_N(_06621_),
    .A2_N(_06635_),
    .B1(_06860_),
    .B2(_06861_),
    .X(_06871_));
 sky130_fd_sc_hd__nand2_1 _29416_ (.A(_06870_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__o211ai_4 _29417_ (.A1(_06683_),
    .A2(_06868_),
    .B1(_06869_),
    .C1(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__a22oi_4 _29418_ (.A1(_06687_),
    .A2(_06837_),
    .B1(_06867_),
    .B2(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__o2bb2ai_1 _29419_ (.A1_N(_06871_),
    .A2_N(_06870_),
    .B1(_06683_),
    .B2(_06868_),
    .Y(_06875_));
 sky130_fd_sc_hd__o21ai_2 _29420_ (.A1(_06685_),
    .A2(_06681_),
    .B1(_06688_),
    .Y(_06876_));
 sky130_fd_sc_hd__o211a_4 _29421_ (.A1(_06866_),
    .A2(_06875_),
    .B1(_06876_),
    .C1(_06867_),
    .X(_06877_));
 sky130_fd_sc_hd__o22ai_4 _29422_ (.A1(_06833_),
    .A2(_06836_),
    .B1(_06874_),
    .B2(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__a21o_1 _29423_ (.A1(_06867_),
    .A2(_06873_),
    .B1(_06876_),
    .X(_06879_));
 sky130_fd_sc_hd__nor2_8 _29424_ (.A(_06836_),
    .B(_06833_),
    .Y(_06880_));
 sky130_fd_sc_hd__nand3_2 _29425_ (.A(_06867_),
    .B(_06876_),
    .C(_06873_),
    .Y(_06881_));
 sky130_fd_sc_hd__nand3_2 _29426_ (.A(_06879_),
    .B(_06880_),
    .C(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__nand3_4 _29427_ (.A(_06878_),
    .B(_06882_),
    .C(_06765_),
    .Y(_06883_));
 sky130_fd_sc_hd__o21ai_2 _29428_ (.A1(_06874_),
    .A2(_06877_),
    .B1(_06880_),
    .Y(_06884_));
 sky130_fd_sc_hd__a21o_1 _29429_ (.A1(_06832_),
    .A2(_06828_),
    .B1(_06835_),
    .X(_06885_));
 sky130_fd_sc_hd__nand3_1 _29430_ (.A(_06832_),
    .B(_06828_),
    .C(_06835_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand2_1 _29431_ (.A(_06885_),
    .B(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__nand3_2 _29432_ (.A(_06879_),
    .B(_06881_),
    .C(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__nand3_4 _29433_ (.A(_06884_),
    .B(_06655_),
    .C(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__nor2_2 _29434_ (.A(_06740_),
    .B(_06693_),
    .Y(_06890_));
 sky130_fd_sc_hd__o2bb2ai_4 _29435_ (.A1_N(_06883_),
    .A2_N(_06889_),
    .B1(_06691_),
    .B2(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_2 _29436_ (.A(_06752_),
    .B(_06745_),
    .Y(_06892_));
 sky130_fd_sc_hd__nand3_4 _29437_ (.A(_06889_),
    .B(_06883_),
    .C(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__clkbuf_4 _29438_ (.A(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__buf_8 _29439_ (.A(_06606_),
    .X(_06895_));
 sky130_fd_sc_hd__a22oi_4 _29440_ (.A1(_06363_),
    .A2(_05451_),
    .B1(_06895_),
    .B2(_05244_),
    .Y(_06896_));
 sky130_fd_sc_hd__nand2_2 _29441_ (.A(_19892_),
    .B(_05456_),
    .Y(_06897_));
 sky130_fd_sc_hd__buf_4 _29442_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06898_));
 sky130_fd_sc_hd__nand2_1 _29443_ (.A(_06898_),
    .B(_05460_),
    .Y(_06899_));
 sky130_fd_sc_hd__nor2_2 _29444_ (.A(_06897_),
    .B(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_2 _29445_ (.A(_06366_),
    .B(_05388_),
    .Y(_06901_));
 sky130_fd_sc_hd__o21bai_2 _29446_ (.A1(_06896_),
    .A2(_06900_),
    .B1_N(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__nand3b_4 _29447_ (.A_N(_06897_),
    .B(_06359_),
    .C(_06199_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_2 _29448_ (.A(_06897_),
    .B(_06899_),
    .Y(_06904_));
 sky130_fd_sc_hd__nand3_4 _29449_ (.A(_06903_),
    .B(_06901_),
    .C(_06904_),
    .Y(_06905_));
 sky130_vsdinv _29450_ (.A(_06612_),
    .Y(_06906_));
 sky130_fd_sc_hd__a21oi_4 _29451_ (.A1(_06906_),
    .A2(_06616_),
    .B1(_06611_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand3_4 _29452_ (.A(_06902_),
    .B(_06905_),
    .C(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__buf_6 _29453_ (.A(_05656_),
    .X(_06909_));
 sky130_fd_sc_hd__a22oi_4 _29454_ (.A1(_06344_),
    .A2(_06249_),
    .B1(_06909_),
    .B2(_20156_),
    .Y(_06910_));
 sky130_fd_sc_hd__nand2_2 _29455_ (.A(_06117_),
    .B(_05664_),
    .Y(_06911_));
 sky130_fd_sc_hd__nand2_2 _29456_ (.A(_06106_),
    .B(_05472_),
    .Y(_06912_));
 sky130_fd_sc_hd__nor2_1 _29457_ (.A(_06911_),
    .B(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__nand2_2 _29458_ (.A(_06051_),
    .B(_05454_),
    .Y(_06914_));
 sky130_fd_sc_hd__o21bai_1 _29459_ (.A1(_06910_),
    .A2(_06913_),
    .B1_N(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand3b_4 _29460_ (.A_N(_06911_),
    .B(_06045_),
    .C(_06473_),
    .Y(_06916_));
 sky130_fd_sc_hd__nand2_1 _29461_ (.A(_06911_),
    .B(_06912_),
    .Y(_06917_));
 sky130_fd_sc_hd__nand3_1 _29462_ (.A(_06916_),
    .B(_06914_),
    .C(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__nand2_2 _29463_ (.A(_06915_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__nand2_2 _29464_ (.A(_06908_),
    .B(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__a21o_2 _29465_ (.A1(_06902_),
    .A2(_06905_),
    .B1(_06907_),
    .X(_06921_));
 sky130_fd_sc_hd__or2b_2 _29466_ (.A(_06920_),
    .B_N(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__a21o_1 _29467_ (.A1(_06921_),
    .A2(_06908_),
    .B1(_06919_),
    .X(_06923_));
 sky130_fd_sc_hd__nor2_2 _29468_ (.A(_06528_),
    .B(_05126_),
    .Y(_06924_));
 sky130_fd_sc_hd__buf_6 _29469_ (.A(_19885_),
    .X(_06925_));
 sky130_fd_sc_hd__nand2_1 _29470_ (.A(_06925_),
    .B(_20173_),
    .Y(_06926_));
 sky130_fd_sc_hd__buf_4 _29471_ (.A(\pcpi_mul.rs2[17] ),
    .X(_06927_));
 sky130_fd_sc_hd__nand2_2 _29472_ (.A(_06927_),
    .B(_20176_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _29473_ (.A(_06926_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__nand2_1 _29474_ (.A(_06924_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__or2_1 _29475_ (.A(_06926_),
    .B(_06928_),
    .X(_06931_));
 sky130_fd_sc_hd__or2b_2 _29476_ (.A(_06930_),
    .B_N(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__a21o_1 _29477_ (.A1(_06931_),
    .A2(_06929_),
    .B1(_06924_),
    .X(_06933_));
 sky130_fd_sc_hd__nand2_4 _29478_ (.A(_06932_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__nand2_1 _29479_ (.A(_06934_),
    .B(_06643_),
    .Y(_06935_));
 sky130_fd_sc_hd__nand3_1 _29480_ (.A(_06932_),
    .B(_06933_),
    .C(_06644_),
    .Y(_06936_));
 sky130_fd_sc_hd__nand2_2 _29481_ (.A(_06935_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__a21o_1 _29482_ (.A1(_06922_),
    .A2(_06923_),
    .B1(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__nand3_4 _29483_ (.A(_06937_),
    .B(_06922_),
    .C(_06923_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand2_4 _29484_ (.A(_06938_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nor2_8 _29485_ (.A(_06940_),
    .B(_06652_),
    .Y(_06941_));
 sky130_fd_sc_hd__and2_2 _29486_ (.A(_06652_),
    .B(_06940_),
    .X(_06942_));
 sky130_fd_sc_hd__nor2_8 _29487_ (.A(_06941_),
    .B(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__a21oi_4 _29488_ (.A1(_06891_),
    .A2(_06894_),
    .B1(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__a21oi_4 _29489_ (.A1(_06889_),
    .A2(_06883_),
    .B1(_06892_),
    .Y(_06945_));
 sky130_fd_sc_hd__nand2_4 _29490_ (.A(_06893_),
    .B(_06943_),
    .Y(_06946_));
 sky130_fd_sc_hd__o21ai_2 _29491_ (.A1(_06945_),
    .A2(_06946_),
    .B1(_06758_),
    .Y(_06947_));
 sky130_fd_sc_hd__nor2_4 _29492_ (.A(_06944_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__o2bb2ai_4 _29493_ (.A1_N(_06894_),
    .A2_N(_06891_),
    .B1(_06941_),
    .B2(_06942_),
    .Y(_06949_));
 sky130_fd_sc_hd__nand3_4 _29494_ (.A(_06891_),
    .B(_06943_),
    .C(_06894_),
    .Y(_06950_));
 sky130_fd_sc_hd__a21oi_4 _29495_ (.A1(_06949_),
    .A2(_06950_),
    .B1(_06758_),
    .Y(_06951_));
 sky130_fd_sc_hd__o22ai_4 _29496_ (.A1(_06794_),
    .A2(_06795_),
    .B1(_06948_),
    .B2(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand2_1 _29497_ (.A(_06748_),
    .B(_06762_),
    .Y(_06953_));
 sky130_fd_sc_hd__nor2_8 _29498_ (.A(_06945_),
    .B(_06946_),
    .Y(_06954_));
 sky130_fd_sc_hd__o22ai_4 _29499_ (.A1(_06761_),
    .A2(_06953_),
    .B1(_06954_),
    .B2(_06944_),
    .Y(_06955_));
 sky130_fd_sc_hd__nand3_4 _29500_ (.A(_06949_),
    .B(_06758_),
    .C(_06950_),
    .Y(_06956_));
 sky130_fd_sc_hd__nor2_4 _29501_ (.A(_06794_),
    .B(_06795_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand3_2 _29502_ (.A(_06955_),
    .B(_06956_),
    .C(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__nand2_1 _29503_ (.A(_06759_),
    .B(_06605_),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_2 _29504_ (.A(_06959_),
    .B(_06768_),
    .Y(_06960_));
 sky130_fd_sc_hd__nand3_4 _29505_ (.A(_06952_),
    .B(_06958_),
    .C(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__o21ai_2 _29506_ (.A1(_06948_),
    .A2(_06951_),
    .B1(_06957_),
    .Y(_06962_));
 sky130_vsdinv _29507_ (.A(_06960_),
    .Y(_06963_));
 sky130_vsdinv _29508_ (.A(_06957_),
    .Y(_06964_));
 sky130_fd_sc_hd__nand3_2 _29509_ (.A(_06955_),
    .B(_06956_),
    .C(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__nand3_4 _29510_ (.A(_06962_),
    .B(_06963_),
    .C(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__o2bb2ai_4 _29511_ (.A1_N(_06961_),
    .A2_N(_06966_),
    .B1(_06576_),
    .B2(_06602_),
    .Y(_06967_));
 sky130_fd_sc_hd__nand2_4 _29512_ (.A(_06966_),
    .B(_06603_),
    .Y(_06968_));
 sky130_fd_sc_hd__nand2_4 _29513_ (.A(_06786_),
    .B(_06779_),
    .Y(_06969_));
 sky130_fd_sc_hd__a21oi_4 _29514_ (.A1(_06967_),
    .A2(_06968_),
    .B1(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__nand3_4 _29515_ (.A(_06967_),
    .B(_06969_),
    .C(_06968_),
    .Y(_06971_));
 sky130_fd_sc_hd__or2b_1 _29516_ (.A(_06970_),
    .B_N(_06971_),
    .X(_06972_));
 sky130_vsdinv _29517_ (.A(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__nand2_1 _29518_ (.A(_06791_),
    .B(_06787_),
    .Y(_06974_));
 sky130_fd_sc_hd__xor2_1 _29519_ (.A(_06973_),
    .B(_06974_),
    .X(_02636_));
 sky130_fd_sc_hd__nand2_1 _29520_ (.A(_06792_),
    .B(_06973_),
    .Y(_06975_));
 sky130_fd_sc_hd__buf_4 _29521_ (.A(_20122_),
    .X(_06976_));
 sky130_fd_sc_hd__nand2_1 _29522_ (.A(_05173_),
    .B(_06816_),
    .Y(_06977_));
 sky130_fd_sc_hd__a21o_1 _29523_ (.A1(_05242_),
    .A2(_06976_),
    .B1(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__buf_4 _29524_ (.A(\pcpi_mul.rs1[17] ),
    .X(_06979_));
 sky130_fd_sc_hd__nand2_1 _29525_ (.A(_05570_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__a21o_1 _29526_ (.A1(_19931_),
    .A2(_20126_),
    .B1(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__nand2_2 _29527_ (.A(_05692_),
    .B(_20130_),
    .Y(_06982_));
 sky130_fd_sc_hd__a21oi_4 _29528_ (.A1(_06978_),
    .A2(_06981_),
    .B1(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__and3_2 _29529_ (.A(_06978_),
    .B(_06981_),
    .C(_06982_),
    .X(_06984_));
 sky130_fd_sc_hd__nor2_2 _29530_ (.A(_06983_),
    .B(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__buf_6 _29531_ (.A(_05227_),
    .X(_06986_));
 sky130_fd_sc_hd__nand2_2 _29532_ (.A(_06986_),
    .B(_06311_),
    .Y(_06987_));
 sky130_fd_sc_hd__buf_6 _29533_ (.A(_19923_),
    .X(_06988_));
 sky130_fd_sc_hd__buf_4 _29534_ (.A(_06293_),
    .X(_06989_));
 sky130_fd_sc_hd__nand2_4 _29535_ (.A(_06988_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__or2_1 _29536_ (.A(_06987_),
    .B(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__nand2_2 _29537_ (.A(_06987_),
    .B(_06990_),
    .Y(_06992_));
 sky130_fd_sc_hd__buf_6 _29538_ (.A(_20117_),
    .X(_06993_));
 sky130_fd_sc_hd__nand2_8 _29539_ (.A(net469),
    .B(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__nand3_2 _29540_ (.A(_06991_),
    .B(_06992_),
    .C(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__a21oi_2 _29541_ (.A1(_06809_),
    .A2(_06803_),
    .B1(_06808_),
    .Y(_06996_));
 sky130_fd_sc_hd__a22oi_4 _29542_ (.A1(_05797_),
    .A2(_20135_),
    .B1(_19925_),
    .B2(_20133_),
    .Y(_06997_));
 sky130_fd_sc_hd__nor2_4 _29543_ (.A(_06987_),
    .B(_06990_),
    .Y(_06998_));
 sky130_vsdinv _29544_ (.A(_06994_),
    .Y(_06999_));
 sky130_fd_sc_hd__o21ai_2 _29545_ (.A1(_06997_),
    .A2(_06998_),
    .B1(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand3_4 _29546_ (.A(_06995_),
    .B(_06996_),
    .C(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__nand2_2 _29547_ (.A(_06802_),
    .B(_06822_),
    .Y(_07002_));
 sky130_fd_sc_hd__buf_6 _29548_ (.A(_06294_),
    .X(_07003_));
 sky130_fd_sc_hd__buf_6 _29549_ (.A(_06311_),
    .X(_07004_));
 sky130_fd_sc_hd__a41oi_4 _29550_ (.A1(_05816_),
    .A2(_05674_),
    .A3(_07003_),
    .A4(_07004_),
    .B1(_06994_),
    .Y(_07005_));
 sky130_fd_sc_hd__nand2_2 _29551_ (.A(_07005_),
    .B(_06992_),
    .Y(_07006_));
 sky130_fd_sc_hd__o21ai_2 _29552_ (.A1(_06997_),
    .A2(_06998_),
    .B1(_06994_),
    .Y(_07007_));
 sky130_fd_sc_hd__nand3_4 _29553_ (.A(_07002_),
    .B(_07006_),
    .C(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__nand3_4 _29554_ (.A(_06985_),
    .B(_07001_),
    .C(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__o2bb2ai_4 _29555_ (.A1_N(_07008_),
    .A2_N(_07001_),
    .B1(_06984_),
    .B2(_06983_),
    .Y(_07010_));
 sky130_vsdinv _29556_ (.A(_06811_),
    .Y(_07011_));
 sky130_fd_sc_hd__o21a_1 _29557_ (.A1(_06820_),
    .A2(_06819_),
    .B1(_06825_),
    .X(_07012_));
 sky130_fd_sc_hd__o2bb2ai_4 _29558_ (.A1_N(_07009_),
    .A2_N(_07010_),
    .B1(_07011_),
    .B2(_07012_),
    .Y(_07013_));
 sky130_vsdinv _29559_ (.A(_06819_),
    .Y(_07014_));
 sky130_fd_sc_hd__o21a_2 _29560_ (.A1(_06815_),
    .A2(_06812_),
    .B1(_07014_),
    .X(_07015_));
 sky130_vsdinv _29561_ (.A(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__nand2_1 _29562_ (.A(_06811_),
    .B(_06821_),
    .Y(_07017_));
 sky130_fd_sc_hd__nand2_1 _29563_ (.A(_07017_),
    .B(_06825_),
    .Y(_07018_));
 sky130_fd_sc_hd__nand3_4 _29564_ (.A(_07018_),
    .B(_07010_),
    .C(_07009_),
    .Y(_07019_));
 sky130_fd_sc_hd__and3_2 _29565_ (.A(_07013_),
    .B(_07016_),
    .C(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__a21oi_4 _29566_ (.A1(_07013_),
    .A2(_07019_),
    .B1(_07016_),
    .Y(_07021_));
 sky130_vsdinv _29567_ (.A(_06855_),
    .Y(_07022_));
 sky130_fd_sc_hd__nor2_2 _29568_ (.A(_06858_),
    .B(_06864_),
    .Y(_07023_));
 sky130_fd_sc_hd__buf_6 _29569_ (.A(_20141_),
    .X(_07024_));
 sky130_fd_sc_hd__a22oi_4 _29570_ (.A1(net468),
    .A2(_05826_),
    .B1(_05499_),
    .B2(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__nand3_4 _29571_ (.A(_06659_),
    .B(_06110_),
    .C(_05822_),
    .Y(_07026_));
 sky130_fd_sc_hd__nor2_4 _29572_ (.A(_05812_),
    .B(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__buf_4 _29573_ (.A(\pcpi_mul.rs1[12] ),
    .X(_07028_));
 sky130_fd_sc_hd__nand2_2 _29574_ (.A(_05601_),
    .B(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__o21ai_2 _29575_ (.A1(_07025_),
    .A2(_07027_),
    .B1(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__o21ai_2 _29576_ (.A1(_06914_),
    .A2(_06910_),
    .B1(_06916_),
    .Y(_07031_));
 sky130_vsdinv _29577_ (.A(_07029_),
    .Y(_07032_));
 sky130_fd_sc_hd__clkbuf_8 _29578_ (.A(_05825_),
    .X(_07033_));
 sky130_fd_sc_hd__a22o_2 _29579_ (.A1(_06478_),
    .A2(_07033_),
    .B1(_06097_),
    .B2(_20142_),
    .X(_07034_));
 sky130_fd_sc_hd__o211ai_4 _29580_ (.A1(_06307_),
    .A2(_07026_),
    .B1(_07032_),
    .C1(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__nand3_4 _29581_ (.A(_07030_),
    .B(_07031_),
    .C(_07035_),
    .Y(_07036_));
 sky130_fd_sc_hd__o21ai_2 _29582_ (.A1(_07025_),
    .A2(_07027_),
    .B1(_07032_),
    .Y(_07037_));
 sky130_fd_sc_hd__o21ai_1 _29583_ (.A1(_06911_),
    .A2(_06912_),
    .B1(_06914_),
    .Y(_07038_));
 sky130_fd_sc_hd__nand2_1 _29584_ (.A(_07038_),
    .B(_06917_),
    .Y(_07039_));
 sky130_fd_sc_hd__o211ai_2 _29585_ (.A1(_06307_),
    .A2(_07026_),
    .B1(_07029_),
    .C1(_07034_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand3_4 _29586_ (.A(_07037_),
    .B(_07039_),
    .C(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__nor2_4 _29587_ (.A(_06847_),
    .B(_06844_),
    .Y(_07042_));
 sky130_fd_sc_hd__o2bb2ai_4 _29588_ (.A1_N(_07036_),
    .A2_N(_07041_),
    .B1(_06842_),
    .B2(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__nor2_2 _29589_ (.A(_06842_),
    .B(_07042_),
    .Y(_07044_));
 sky130_fd_sc_hd__nand3_4 _29590_ (.A(_07036_),
    .B(_07041_),
    .C(_07044_),
    .Y(_07045_));
 sky130_fd_sc_hd__nand2_4 _29591_ (.A(_06920_),
    .B(_06921_),
    .Y(_07046_));
 sky130_fd_sc_hd__a21oi_4 _29592_ (.A1(_07043_),
    .A2(_07045_),
    .B1(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__and3_1 _29593_ (.A(_07030_),
    .B(_07031_),
    .C(_07035_),
    .X(_07048_));
 sky130_fd_sc_hd__nand2_1 _29594_ (.A(_07041_),
    .B(_07044_),
    .Y(_07049_));
 sky130_fd_sc_hd__o211a_1 _29595_ (.A1(_07048_),
    .A2(_07049_),
    .B1(_07043_),
    .C1(_07046_),
    .X(_07050_));
 sky130_fd_sc_hd__o22ai_4 _29596_ (.A1(_07022_),
    .A2(_07023_),
    .B1(_07047_),
    .B2(_07050_),
    .Y(_07051_));
 sky130_vsdinv _29597_ (.A(_06859_),
    .Y(_07052_));
 sky130_fd_sc_hd__nand3_4 _29598_ (.A(_07046_),
    .B(_07043_),
    .C(_07045_),
    .Y(_07053_));
 sky130_fd_sc_hd__nand2_1 _29599_ (.A(_07043_),
    .B(_07045_),
    .Y(_07054_));
 sky130_fd_sc_hd__and2_1 _29600_ (.A(_06920_),
    .B(_06921_),
    .X(_07055_));
 sky130_fd_sc_hd__nand2_2 _29601_ (.A(_07054_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__o211ai_4 _29602_ (.A1(_06864_),
    .A2(_07052_),
    .B1(_07053_),
    .C1(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__and2_1 _29603_ (.A(_06682_),
    .B(_06668_),
    .X(_07058_));
 sky130_fd_sc_hd__o21ai_4 _29604_ (.A1(_07058_),
    .A2(_06863_),
    .B1(_06869_),
    .Y(_07059_));
 sky130_fd_sc_hd__a21oi_4 _29605_ (.A1(_07051_),
    .A2(_07057_),
    .B1(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__o2bb2ai_1 _29606_ (.A1_N(_07055_),
    .A2_N(_07054_),
    .B1(_06864_),
    .B2(_07052_),
    .Y(_07061_));
 sky130_fd_sc_hd__o211a_2 _29607_ (.A1(_07050_),
    .A2(_07061_),
    .B1(_07059_),
    .C1(_07051_),
    .X(_07062_));
 sky130_fd_sc_hd__o22ai_4 _29608_ (.A1(_07020_),
    .A2(_07021_),
    .B1(_07060_),
    .B2(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__a21o_1 _29609_ (.A1(_07051_),
    .A2(_07057_),
    .B1(_07059_),
    .X(_07064_));
 sky130_fd_sc_hd__nor2_4 _29610_ (.A(_07021_),
    .B(_07020_),
    .Y(_07065_));
 sky130_fd_sc_hd__nand3_4 _29611_ (.A(_07051_),
    .B(_07059_),
    .C(_07057_),
    .Y(_07066_));
 sky130_fd_sc_hd__nand3_2 _29612_ (.A(_07064_),
    .B(_07065_),
    .C(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__nand3_4 _29613_ (.A(_07063_),
    .B(_07067_),
    .C(_06941_),
    .Y(_07068_));
 sky130_fd_sc_hd__o21ai_2 _29614_ (.A1(_07060_),
    .A2(_07062_),
    .B1(_07065_),
    .Y(_07069_));
 sky130_vsdinv _29615_ (.A(_06941_),
    .Y(_07070_));
 sky130_fd_sc_hd__a21o_1 _29616_ (.A1(_07013_),
    .A2(_07019_),
    .B1(_07016_),
    .X(_07071_));
 sky130_fd_sc_hd__nand3_1 _29617_ (.A(_07013_),
    .B(_07016_),
    .C(_07019_),
    .Y(_07072_));
 sky130_fd_sc_hd__nand2_2 _29618_ (.A(_07071_),
    .B(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__nand3_2 _29619_ (.A(_07064_),
    .B(_07066_),
    .C(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__nand3_4 _29620_ (.A(_07069_),
    .B(_07070_),
    .C(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__nor2_8 _29621_ (.A(_06877_),
    .B(_06880_),
    .Y(_07076_));
 sky130_fd_sc_hd__o2bb2ai_2 _29622_ (.A1_N(_07068_),
    .A2_N(_07075_),
    .B1(_06874_),
    .B2(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__nor2_1 _29623_ (.A(_06926_),
    .B(_06928_),
    .Y(_07078_));
 sky130_fd_sc_hd__o211a_1 _29624_ (.A1(_07078_),
    .A2(_06930_),
    .B1(_06643_),
    .C1(_06933_),
    .X(_07079_));
 sky130_fd_sc_hd__nand2_4 _29625_ (.A(_06927_),
    .B(_20173_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand2_4 _29626_ (.A(_06925_),
    .B(_20170_),
    .Y(_07081_));
 sky130_fd_sc_hd__nor2_8 _29627_ (.A(_07080_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__nand2_2 _29628_ (.A(_06640_),
    .B(_06551_),
    .Y(_07083_));
 sky130_vsdinv _29629_ (.A(_07083_),
    .Y(_07084_));
 sky130_fd_sc_hd__nand2_2 _29630_ (.A(_07080_),
    .B(_07081_),
    .Y(_07085_));
 sky130_fd_sc_hd__nand2_2 _29631_ (.A(_07084_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__clkbuf_4 _29632_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07087_));
 sky130_fd_sc_hd__buf_6 _29633_ (.A(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__clkbuf_4 _29634_ (.A(_19885_),
    .X(_07089_));
 sky130_fd_sc_hd__buf_6 _29635_ (.A(_07089_),
    .X(_07090_));
 sky130_fd_sc_hd__a22oi_4 _29636_ (.A1(_07088_),
    .A2(_05146_),
    .B1(_07090_),
    .B2(_20171_),
    .Y(_07091_));
 sky130_fd_sc_hd__o21ai_2 _29637_ (.A1(_07091_),
    .A2(_07082_),
    .B1(_07083_),
    .Y(_07092_));
 sky130_fd_sc_hd__o21ai_1 _29638_ (.A1(_07082_),
    .A2(_07086_),
    .B1(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__a21oi_1 _29639_ (.A1(_06924_),
    .A2(_06929_),
    .B1(_07078_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2_2 _29640_ (.A(_07093_),
    .B(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__nand2_1 _29641_ (.A(_06930_),
    .B(_06931_),
    .Y(_07096_));
 sky130_fd_sc_hd__o211ai_4 _29642_ (.A1(_07082_),
    .A2(_07086_),
    .B1(_07092_),
    .C1(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__nand3_4 _29643_ (.A(_07079_),
    .B(_07095_),
    .C(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__nand2_2 _29644_ (.A(_07095_),
    .B(_07097_),
    .Y(_07099_));
 sky130_fd_sc_hd__o21ai_4 _29645_ (.A1(_06644_),
    .A2(_06934_),
    .B1(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__nand2_1 _29646_ (.A(_07098_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__clkbuf_8 _29647_ (.A(\pcpi_mul.rs2[14] ),
    .X(_07102_));
 sky130_fd_sc_hd__nand2_4 _29648_ (.A(_07102_),
    .B(_05237_),
    .Y(_07103_));
 sky130_fd_sc_hd__nand2_4 _29649_ (.A(_06898_),
    .B(_05289_),
    .Y(_07104_));
 sky130_fd_sc_hd__nor2_8 _29650_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__nand2_2 _29651_ (.A(_19898_),
    .B(_20158_),
    .Y(_07106_));
 sky130_vsdinv _29652_ (.A(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__nand2_2 _29653_ (.A(_07103_),
    .B(_07104_),
    .Y(_07108_));
 sky130_fd_sc_hd__nand2_2 _29654_ (.A(_07107_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__o21ai_2 _29655_ (.A1(_06901_),
    .A2(_06896_),
    .B1(_06903_),
    .Y(_07110_));
 sky130_fd_sc_hd__a22oi_4 _29656_ (.A1(_06544_),
    .A2(_20165_),
    .B1(_06546_),
    .B2(_05481_),
    .Y(_07111_));
 sky130_fd_sc_hd__o21ai_2 _29657_ (.A1(_07111_),
    .A2(_07105_),
    .B1(_07106_),
    .Y(_07112_));
 sky130_fd_sc_hd__o211ai_4 _29658_ (.A1(_07105_),
    .A2(_07109_),
    .B1(_07110_),
    .C1(_07112_),
    .Y(_07113_));
 sky130_fd_sc_hd__o21ai_2 _29659_ (.A1(_07111_),
    .A2(_07105_),
    .B1(_07107_),
    .Y(_07114_));
 sky130_fd_sc_hd__buf_6 _29660_ (.A(_19895_),
    .X(_07115_));
 sky130_fd_sc_hd__nand3b_2 _29661_ (.A_N(_07103_),
    .B(_07115_),
    .C(_06348_),
    .Y(_07116_));
 sky130_fd_sc_hd__nand3_2 _29662_ (.A(_07116_),
    .B(_07106_),
    .C(_07108_),
    .Y(_07117_));
 sky130_vsdinv _29663_ (.A(_06901_),
    .Y(_07118_));
 sky130_fd_sc_hd__a21oi_2 _29664_ (.A1(_07118_),
    .A2(_06904_),
    .B1(_06900_),
    .Y(_07119_));
 sky130_fd_sc_hd__nand3_4 _29665_ (.A(_07114_),
    .B(_07117_),
    .C(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__a22oi_4 _29666_ (.A1(_06531_),
    .A2(_06473_),
    .B1(_06196_),
    .B2(_06476_),
    .Y(_07121_));
 sky130_fd_sc_hd__nand2_1 _29667_ (.A(_06041_),
    .B(_06472_),
    .Y(_07122_));
 sky130_fd_sc_hd__nand2_1 _29668_ (.A(_06631_),
    .B(_05831_),
    .Y(_07123_));
 sky130_fd_sc_hd__nor2_1 _29669_ (.A(_07122_),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__nand2_2 _29670_ (.A(_05952_),
    .B(_20149_),
    .Y(_07125_));
 sky130_vsdinv _29671_ (.A(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__o21ai_1 _29672_ (.A1(_07121_),
    .A2(_07124_),
    .B1(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand3b_2 _29673_ (.A_N(_07122_),
    .B(_06107_),
    .C(_05979_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand2_1 _29674_ (.A(_07122_),
    .B(_07123_),
    .Y(_07129_));
 sky130_fd_sc_hd__nand3_1 _29675_ (.A(_07128_),
    .B(_07129_),
    .C(_07125_),
    .Y(_07130_));
 sky130_fd_sc_hd__nand2_2 _29676_ (.A(_07127_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__a21o_1 _29677_ (.A1(_07113_),
    .A2(_07120_),
    .B1(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand3_4 _29678_ (.A(_07113_),
    .B(_07120_),
    .C(_07131_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_2 _29679_ (.A(_07132_),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nand2_1 _29680_ (.A(_07101_),
    .B(_07134_),
    .Y(_07135_));
 sky130_fd_sc_hd__nand3b_4 _29681_ (.A_N(_07134_),
    .B(_07100_),
    .C(_07098_),
    .Y(_07136_));
 sky130_fd_sc_hd__nand3b_4 _29682_ (.A_N(_06939_),
    .B(_07135_),
    .C(_07136_),
    .Y(_07137_));
 sky130_fd_sc_hd__a21o_1 _29683_ (.A1(_07098_),
    .A2(_07100_),
    .B1(_07134_),
    .X(_07138_));
 sky130_fd_sc_hd__nand3_2 _29684_ (.A(_07134_),
    .B(_07098_),
    .C(_07100_),
    .Y(_07139_));
 sky130_fd_sc_hd__nand3_4 _29685_ (.A(_07138_),
    .B(_06939_),
    .C(_07139_),
    .Y(_07140_));
 sky130_vsdinv _29686_ (.A(_19877_),
    .Y(_07141_));
 sky130_fd_sc_hd__nor2_8 _29687_ (.A(_07141_),
    .B(_04841_),
    .Y(_07142_));
 sky130_fd_sc_hd__a21oi_4 _29688_ (.A1(_07137_),
    .A2(_07140_),
    .B1(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__and3_4 _29689_ (.A(_07137_),
    .B(_07140_),
    .C(_07142_),
    .X(_07144_));
 sky130_fd_sc_hd__nor2_4 _29690_ (.A(_07143_),
    .B(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__nor2_4 _29691_ (.A(_06874_),
    .B(_07076_),
    .Y(_07146_));
 sky130_fd_sc_hd__nand3_4 _29692_ (.A(_07075_),
    .B(_07146_),
    .C(_07068_),
    .Y(_07147_));
 sky130_fd_sc_hd__nand3_4 _29693_ (.A(_07077_),
    .B(_07145_),
    .C(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__buf_2 _29694_ (.A(_07068_),
    .X(_07149_));
 sky130_fd_sc_hd__a2bb2oi_4 _29695_ (.A1_N(_06874_),
    .A2_N(_07076_),
    .B1(_07149_),
    .B2(_07075_),
    .Y(_07150_));
 sky130_fd_sc_hd__nor2_1 _29696_ (.A(_06874_),
    .B(_06887_),
    .Y(_07151_));
 sky130_fd_sc_hd__o211a_1 _29697_ (.A1(_06877_),
    .A2(_07151_),
    .B1(_07149_),
    .C1(_07075_),
    .X(_07152_));
 sky130_fd_sc_hd__o22ai_4 _29698_ (.A1(_07144_),
    .A2(_07143_),
    .B1(_07150_),
    .B2(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__a2bb2oi_4 _29699_ (.A1_N(_06945_),
    .A2_N(_06946_),
    .B1(_07148_),
    .B2(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__nand2_2 _29700_ (.A(_07147_),
    .B(_07145_),
    .Y(_07155_));
 sky130_fd_sc_hd__o211a_1 _29701_ (.A1(_07150_),
    .A2(_07155_),
    .B1(_06954_),
    .C1(_07153_),
    .X(_07156_));
 sky130_vsdinv _29702_ (.A(_06832_),
    .Y(_07157_));
 sky130_fd_sc_hd__o21a_2 _29703_ (.A1(_06834_),
    .A2(_07157_),
    .B1(_06828_),
    .X(_07158_));
 sky130_fd_sc_hd__a21o_2 _29704_ (.A1(_06894_),
    .A2(_06883_),
    .B1(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__nand3_2 _29705_ (.A(_06894_),
    .B(_06883_),
    .C(_07158_),
    .Y(_07160_));
 sky130_fd_sc_hd__nand2_4 _29706_ (.A(_07159_),
    .B(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__o21bai_2 _29707_ (.A1(_07154_),
    .A2(_07156_),
    .B1_N(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__a21oi_2 _29708_ (.A1(_06955_),
    .A2(_06957_),
    .B1(_06948_),
    .Y(_07163_));
 sky130_fd_sc_hd__a21o_1 _29709_ (.A1(_07153_),
    .A2(_07148_),
    .B1(_06954_),
    .X(_07164_));
 sky130_fd_sc_hd__nand3_4 _29710_ (.A(_07153_),
    .B(_06954_),
    .C(_07148_),
    .Y(_07165_));
 sky130_fd_sc_hd__nand3_2 _29711_ (.A(_07164_),
    .B(_07165_),
    .C(_07161_),
    .Y(_07166_));
 sky130_fd_sc_hd__nand3_4 _29712_ (.A(_07162_),
    .B(_07163_),
    .C(_07166_),
    .Y(_07167_));
 sky130_fd_sc_hd__nand2_4 _29713_ (.A(_07167_),
    .B(_06794_),
    .Y(_07168_));
 sky130_fd_sc_hd__o21ai_2 _29714_ (.A1(_07154_),
    .A2(_07156_),
    .B1(_07161_),
    .Y(_07169_));
 sky130_fd_sc_hd__o21ai_2 _29715_ (.A1(_06964_),
    .A2(_06951_),
    .B1(_06956_),
    .Y(_07170_));
 sky130_fd_sc_hd__nand3b_4 _29716_ (.A_N(_07161_),
    .B(_07164_),
    .C(_07165_),
    .Y(_07171_));
 sky130_fd_sc_hd__nand3_4 _29717_ (.A(_07169_),
    .B(_07170_),
    .C(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__nand2_1 _29718_ (.A(_07172_),
    .B(_07167_),
    .Y(_07173_));
 sky130_vsdinv _29719_ (.A(_06794_),
    .Y(_07174_));
 sky130_fd_sc_hd__a22oi_4 _29720_ (.A1(_06968_),
    .A2(_06961_),
    .B1(_07173_),
    .B2(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__o2bb2ai_2 _29721_ (.A1_N(_07167_),
    .A2_N(_07172_),
    .B1(_06762_),
    .B2(_06793_),
    .Y(_07176_));
 sky130_fd_sc_hd__nand2_1 _29722_ (.A(_06968_),
    .B(_06961_),
    .Y(_07177_));
 sky130_fd_sc_hd__a21oi_2 _29723_ (.A1(_07176_),
    .A2(_07168_),
    .B1(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__a21oi_4 _29724_ (.A1(_07168_),
    .A2(_07175_),
    .B1(_07178_),
    .Y(_07179_));
 sky130_vsdinv _29725_ (.A(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__a21oi_4 _29726_ (.A1(_06787_),
    .A2(_06971_),
    .B1(_06970_),
    .Y(_07181_));
 sky130_vsdinv _29727_ (.A(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__and3_1 _29728_ (.A(_06975_),
    .B(_07180_),
    .C(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__a21o_1 _29729_ (.A1(_06975_),
    .A2(_07182_),
    .B1(_07180_),
    .X(_07184_));
 sky130_fd_sc_hd__nor2b_1 _29730_ (.A(_07183_),
    .B_N(_07184_),
    .Y(_02637_));
 sky130_fd_sc_hd__buf_6 _29731_ (.A(_05985_),
    .X(_07185_));
 sky130_fd_sc_hd__a22oi_4 _29732_ (.A1(_06483_),
    .A2(_05999_),
    .B1(_19915_),
    .B2(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__nand3_4 _29733_ (.A(_19911_),
    .B(_06110_),
    .C(_06153_),
    .Y(_07187_));
 sky130_fd_sc_hd__nor2_8 _29734_ (.A(_06445_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__nand2_2 _29735_ (.A(_05601_),
    .B(_06311_),
    .Y(_07189_));
 sky130_fd_sc_hd__o21ai_2 _29736_ (.A1(_07186_),
    .A2(_07188_),
    .B1(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__clkbuf_8 _29737_ (.A(_06445_),
    .X(_07191_));
 sky130_vsdinv _29738_ (.A(_07189_),
    .Y(_07192_));
 sky130_fd_sc_hd__a22o_1 _29739_ (.A1(_06100_),
    .A2(_06154_),
    .B1(_06474_),
    .B2(_07185_),
    .X(_07193_));
 sky130_fd_sc_hd__o211ai_2 _29740_ (.A1(_07191_),
    .A2(_07187_),
    .B1(_07192_),
    .C1(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__o21ai_2 _29741_ (.A1(_07125_),
    .A2(_07121_),
    .B1(_07128_),
    .Y(_07195_));
 sky130_fd_sc_hd__nand3_4 _29742_ (.A(_07190_),
    .B(_07194_),
    .C(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__o21ai_2 _29743_ (.A1(_07186_),
    .A2(_07188_),
    .B1(_07192_),
    .Y(_07197_));
 sky130_fd_sc_hd__a21oi_2 _29744_ (.A1(_07126_),
    .A2(_07129_),
    .B1(_07124_),
    .Y(_07198_));
 sky130_fd_sc_hd__o211ai_4 _29745_ (.A1(_07191_),
    .A2(_07187_),
    .B1(_07189_),
    .C1(_07193_),
    .Y(_07199_));
 sky130_fd_sc_hd__nand3_4 _29746_ (.A(_07197_),
    .B(_07198_),
    .C(_07199_),
    .Y(_07200_));
 sky130_fd_sc_hd__nor2_4 _29747_ (.A(_07032_),
    .B(_07027_),
    .Y(_07201_));
 sky130_fd_sc_hd__o2bb2ai_4 _29748_ (.A1_N(_07196_),
    .A2_N(_07200_),
    .B1(_07025_),
    .B2(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__nor2_4 _29749_ (.A(_07025_),
    .B(_07201_),
    .Y(_07203_));
 sky130_fd_sc_hd__nand3_4 _29750_ (.A(_07200_),
    .B(_07196_),
    .C(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__nand2_1 _29751_ (.A(_07120_),
    .B(_07131_),
    .Y(_07205_));
 sky130_fd_sc_hd__nand2_4 _29752_ (.A(_07205_),
    .B(_07113_),
    .Y(_07206_));
 sky130_fd_sc_hd__a21oi_4 _29753_ (.A1(_07202_),
    .A2(_07204_),
    .B1(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__nand2_1 _29754_ (.A(_07200_),
    .B(_07203_),
    .Y(_07208_));
 sky130_vsdinv _29755_ (.A(_07196_),
    .Y(_07209_));
 sky130_fd_sc_hd__o211a_1 _29756_ (.A1(_07208_),
    .A2(_07209_),
    .B1(_07202_),
    .C1(_07206_),
    .X(_07210_));
 sky130_fd_sc_hd__nand2_2 _29757_ (.A(_07049_),
    .B(_07036_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21bai_2 _29758_ (.A1(_07207_),
    .A2(_07210_),
    .B1_N(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__and2_1 _29759_ (.A(_06865_),
    .B(_06851_),
    .X(_07213_));
 sky130_fd_sc_hd__o21ai_2 _29760_ (.A1(_07213_),
    .A2(_07047_),
    .B1(_07053_),
    .Y(_07214_));
 sky130_fd_sc_hd__a21o_1 _29761_ (.A1(_07202_),
    .A2(_07204_),
    .B1(_07206_),
    .X(_07215_));
 sky130_fd_sc_hd__nand3_4 _29762_ (.A(_07206_),
    .B(_07202_),
    .C(_07204_),
    .Y(_07216_));
 sky130_fd_sc_hd__nand3_2 _29763_ (.A(_07215_),
    .B(_07216_),
    .C(_07211_),
    .Y(_07217_));
 sky130_fd_sc_hd__nand3_4 _29764_ (.A(_07212_),
    .B(_07214_),
    .C(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__o21ai_2 _29765_ (.A1(_07207_),
    .A2(_07210_),
    .B1(_07211_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_1 _29766_ (.A(_07053_),
    .B(_07213_),
    .Y(_07220_));
 sky130_fd_sc_hd__nand2_1 _29767_ (.A(_07220_),
    .B(_07056_),
    .Y(_07221_));
 sky130_vsdinv _29768_ (.A(_07211_),
    .Y(_07222_));
 sky130_fd_sc_hd__nand3_2 _29769_ (.A(_07215_),
    .B(_07216_),
    .C(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__nand3_4 _29770_ (.A(_07219_),
    .B(_07221_),
    .C(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__a21o_1 _29771_ (.A1(_06978_),
    .A2(_06981_),
    .B1(_06982_),
    .X(_07225_));
 sky130_fd_sc_hd__o21a_4 _29772_ (.A1(_06977_),
    .A2(_06980_),
    .B1(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__a21oi_2 _29773_ (.A1(_07007_),
    .A2(_07006_),
    .B1(_07002_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand3_1 _29774_ (.A(_06978_),
    .B(_06981_),
    .C(_06982_),
    .Y(_07228_));
 sky130_fd_sc_hd__nand2_2 _29775_ (.A(_07225_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__o21a_2 _29776_ (.A1(_07227_),
    .A2(_07229_),
    .B1(_07008_),
    .X(_07230_));
 sky130_fd_sc_hd__a21oi_4 _29777_ (.A1(_06999_),
    .A2(_06992_),
    .B1(_06998_),
    .Y(_07231_));
 sky130_fd_sc_hd__buf_4 _29778_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07232_));
 sky130_fd_sc_hd__buf_6 _29779_ (.A(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__nand2_8 _29780_ (.A(_19937_),
    .B(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__a22oi_4 _29781_ (.A1(_05376_),
    .A2(_06989_),
    .B1(_05377_),
    .B2(_06719_),
    .Y(_07235_));
 sky130_fd_sc_hd__nor2_1 _29782_ (.A(_07234_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__nand2_2 _29783_ (.A(_05311_),
    .B(_06989_),
    .Y(_07237_));
 sky130_fd_sc_hd__nand2_2 _29784_ (.A(_05312_),
    .B(_06719_),
    .Y(_07238_));
 sky130_fd_sc_hd__or2_4 _29785_ (.A(_07237_),
    .B(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__nand2_1 _29786_ (.A(_07236_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__nor2_2 _29787_ (.A(_07237_),
    .B(_07238_),
    .Y(_07241_));
 sky130_fd_sc_hd__o21ai_2 _29788_ (.A1(_07235_),
    .A2(_07241_),
    .B1(_07234_),
    .Y(_07242_));
 sky130_fd_sc_hd__nand3b_4 _29789_ (.A_N(_07231_),
    .B(_07240_),
    .C(_07242_),
    .Y(_07243_));
 sky130_vsdinv _29790_ (.A(_07235_),
    .Y(_07244_));
 sky130_fd_sc_hd__nand3_2 _29791_ (.A(_07239_),
    .B(_07244_),
    .C(_07234_),
    .Y(_07245_));
 sky130_fd_sc_hd__o21bai_2 _29792_ (.A1(_07235_),
    .A2(_07241_),
    .B1_N(_07234_),
    .Y(_07246_));
 sky130_fd_sc_hd__nand3_4 _29793_ (.A(_07245_),
    .B(_07231_),
    .C(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__nand2_1 _29794_ (.A(_07243_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__buf_4 _29795_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07249_));
 sky130_fd_sc_hd__buf_6 _29796_ (.A(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__buf_6 _29797_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07251_));
 sky130_fd_sc_hd__nand2_2 _29798_ (.A(_05139_),
    .B(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__a21o_2 _29799_ (.A1(_05821_),
    .A2(_07250_),
    .B1(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__buf_4 _29800_ (.A(_20117_),
    .X(_07254_));
 sky130_fd_sc_hd__nand2_4 _29801_ (.A(_05141_),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__a21o_2 _29802_ (.A1(_06314_),
    .A2(_06976_),
    .B1(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__buf_6 _29803_ (.A(\pcpi_mul.rs1[16] ),
    .X(_07257_));
 sky130_fd_sc_hd__buf_6 _29804_ (.A(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__nand2_4 _29805_ (.A(_05692_),
    .B(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__a21oi_4 _29806_ (.A1(_07253_),
    .A2(_07256_),
    .B1(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__and3_1 _29807_ (.A(_07253_),
    .B(_07256_),
    .C(_07259_),
    .X(_07261_));
 sky130_fd_sc_hd__nor2_4 _29808_ (.A(_07260_),
    .B(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__nand2_2 _29809_ (.A(_07248_),
    .B(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__nand3_1 _29810_ (.A(_07253_),
    .B(_07256_),
    .C(_07259_),
    .Y(_07264_));
 sky130_fd_sc_hd__or2b_2 _29811_ (.A(_07260_),
    .B_N(_07264_),
    .X(_07265_));
 sky130_fd_sc_hd__nand3_4 _29812_ (.A(_07265_),
    .B(_07247_),
    .C(_07243_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand3_4 _29813_ (.A(_07230_),
    .B(_07263_),
    .C(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_1 _29814_ (.A(_07248_),
    .B(_07265_),
    .Y(_07268_));
 sky130_fd_sc_hd__o21ai_2 _29815_ (.A1(_07227_),
    .A2(_07229_),
    .B1(_07008_),
    .Y(_07269_));
 sky130_fd_sc_hd__nand3_2 _29816_ (.A(_07262_),
    .B(_07247_),
    .C(_07243_),
    .Y(_07270_));
 sky130_fd_sc_hd__nand3_4 _29817_ (.A(_07268_),
    .B(_07269_),
    .C(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_1 _29818_ (.A(_07267_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__nor2_4 _29819_ (.A(_07226_),
    .B(_07272_),
    .Y(_07273_));
 sky130_fd_sc_hd__a21boi_4 _29820_ (.A1(_07267_),
    .A2(_07271_),
    .B1_N(_07226_),
    .Y(_07274_));
 sky130_fd_sc_hd__o2bb2ai_2 _29821_ (.A1_N(_07218_),
    .A2_N(_07224_),
    .B1(_07273_),
    .B2(_07274_),
    .Y(_07275_));
 sky130_vsdinv _29822_ (.A(_07137_),
    .Y(_07276_));
 sky130_fd_sc_hd__a31oi_4 _29823_ (.A1(_07230_),
    .A2(_07263_),
    .A3(_07266_),
    .B1(_07226_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21oi_2 _29824_ (.A1(_07271_),
    .A2(_07277_),
    .B1(_07274_),
    .Y(_07278_));
 sky130_fd_sc_hd__nand3_2 _29825_ (.A(_07278_),
    .B(_07224_),
    .C(_07218_),
    .Y(_07279_));
 sky130_fd_sc_hd__nand3_4 _29826_ (.A(_07275_),
    .B(_07276_),
    .C(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__nand2_1 _29827_ (.A(_07224_),
    .B(_07218_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand2_1 _29828_ (.A(_07281_),
    .B(_07278_),
    .Y(_07282_));
 sky130_fd_sc_hd__o211ai_4 _29829_ (.A1(_07274_),
    .A2(_07273_),
    .B1(_07224_),
    .C1(_07218_),
    .Y(_07283_));
 sky130_fd_sc_hd__nand3_4 _29830_ (.A(_07282_),
    .B(_07137_),
    .C(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__nor2_2 _29831_ (.A(_07062_),
    .B(_07065_),
    .Y(_07285_));
 sky130_fd_sc_hd__o2bb2ai_4 _29832_ (.A1_N(_07280_),
    .A2_N(_07284_),
    .B1(_07060_),
    .B2(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__o21ai_2 _29833_ (.A1(_07073_),
    .A2(_07060_),
    .B1(_07066_),
    .Y(_07287_));
 sky130_fd_sc_hd__nand3_4 _29834_ (.A(_07284_),
    .B(_07280_),
    .C(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__buf_6 _29835_ (.A(_07087_),
    .X(_07289_));
 sky130_fd_sc_hd__nand2_2 _29836_ (.A(_07289_),
    .B(_05300_),
    .Y(_07290_));
 sky130_fd_sc_hd__clkbuf_8 _29837_ (.A(_07089_),
    .X(_07291_));
 sky130_fd_sc_hd__nand2_2 _29838_ (.A(_07291_),
    .B(_20168_),
    .Y(_07292_));
 sky130_fd_sc_hd__or2_2 _29839_ (.A(_07290_),
    .B(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__buf_6 _29840_ (.A(_07087_),
    .X(_07294_));
 sky130_fd_sc_hd__buf_6 _29841_ (.A(_06636_),
    .X(_07295_));
 sky130_fd_sc_hd__a22oi_4 _29842_ (.A1(_07294_),
    .A2(_05143_),
    .B1(_07295_),
    .B2(_05182_),
    .Y(_07296_));
 sky130_vsdinv _29843_ (.A(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__nand2_2 _29844_ (.A(_06640_),
    .B(_05549_),
    .Y(_07298_));
 sky130_fd_sc_hd__nand3_2 _29845_ (.A(_07293_),
    .B(_07297_),
    .C(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__a21oi_4 _29846_ (.A1(_07084_),
    .A2(_07085_),
    .B1(_07082_),
    .Y(_07300_));
 sky130_fd_sc_hd__nor2_4 _29847_ (.A(_07290_),
    .B(_07292_),
    .Y(_07301_));
 sky130_vsdinv _29848_ (.A(_07298_),
    .Y(_07302_));
 sky130_fd_sc_hd__o21ai_2 _29849_ (.A1(_07296_),
    .A2(_07301_),
    .B1(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand3_4 _29850_ (.A(_07299_),
    .B(_07300_),
    .C(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__nand3_2 _29851_ (.A(_07293_),
    .B(_07297_),
    .C(_07302_),
    .Y(_07305_));
 sky130_fd_sc_hd__o21ai_2 _29852_ (.A1(_07296_),
    .A2(_07301_),
    .B1(_07298_),
    .Y(_07306_));
 sky130_fd_sc_hd__nand3b_4 _29853_ (.A_N(_07300_),
    .B(_07305_),
    .C(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__nand3b_4 _29854_ (.A_N(_07097_),
    .B(_07304_),
    .C(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__nand2_1 _29855_ (.A(_07307_),
    .B(_07304_),
    .Y(_07309_));
 sky130_fd_sc_hd__nand2_2 _29856_ (.A(_07309_),
    .B(_07097_),
    .Y(_07310_));
 sky130_fd_sc_hd__nand2_1 _29857_ (.A(_07109_),
    .B(_07116_),
    .Y(_07311_));
 sky130_fd_sc_hd__a22oi_4 _29858_ (.A1(_06357_),
    .A2(_05286_),
    .B1(_06895_),
    .B2(_06249_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand2_2 _29859_ (.A(_06543_),
    .B(_05285_),
    .Y(_07313_));
 sky130_fd_sc_hd__nand2_2 _29860_ (.A(_06898_),
    .B(_05391_),
    .Y(_07314_));
 sky130_fd_sc_hd__nor2_4 _29861_ (.A(_07313_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand2_2 _29862_ (.A(_19898_),
    .B(_06472_),
    .Y(_07316_));
 sky130_fd_sc_hd__o21ai_2 _29863_ (.A1(_07312_),
    .A2(_07315_),
    .B1(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__nand3b_4 _29864_ (.A_N(_07313_),
    .B(_19896_),
    .C(_05474_),
    .Y(_07318_));
 sky130_vsdinv _29865_ (.A(_07316_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand2_2 _29866_ (.A(_07313_),
    .B(_07314_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand3_2 _29867_ (.A(_07318_),
    .B(_07319_),
    .C(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nand3_4 _29868_ (.A(_07311_),
    .B(_07317_),
    .C(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__o21ai_2 _29869_ (.A1(_07312_),
    .A2(_07315_),
    .B1(_07319_),
    .Y(_07323_));
 sky130_fd_sc_hd__nand3_2 _29870_ (.A(_07318_),
    .B(_07316_),
    .C(_07320_),
    .Y(_07324_));
 sky130_fd_sc_hd__a21oi_2 _29871_ (.A1(_07107_),
    .A2(_07108_),
    .B1(_07105_),
    .Y(_07325_));
 sky130_fd_sc_hd__nand3_4 _29872_ (.A(_07323_),
    .B(_07324_),
    .C(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__a22oi_4 _29873_ (.A1(_06118_),
    .A2(_05463_),
    .B1(_05657_),
    .B2(_06289_),
    .Y(_07327_));
 sky130_fd_sc_hd__nand2_1 _29874_ (.A(_06041_),
    .B(_06475_),
    .Y(_07328_));
 sky130_fd_sc_hd__nand2_1 _29875_ (.A(_06106_),
    .B(_05827_),
    .Y(_07329_));
 sky130_fd_sc_hd__nor2_2 _29876_ (.A(_07328_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_2 _29877_ (.A(_05952_),
    .B(_05826_),
    .Y(_07331_));
 sky130_fd_sc_hd__o21bai_2 _29878_ (.A1(_07327_),
    .A2(_07330_),
    .B1_N(_07331_),
    .Y(_07332_));
 sky130_fd_sc_hd__clkbuf_8 _29879_ (.A(_06106_),
    .X(_07333_));
 sky130_fd_sc_hd__nand3b_4 _29880_ (.A_N(_07328_),
    .B(_07333_),
    .C(_05820_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_1 _29881_ (.A(_07328_),
    .B(_07329_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand3_2 _29882_ (.A(_07334_),
    .B(_07331_),
    .C(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__nand2_4 _29883_ (.A(_07332_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__a21oi_1 _29884_ (.A1(_07322_),
    .A2(_07326_),
    .B1(_07337_),
    .Y(_07338_));
 sky130_vsdinv _29885_ (.A(_07337_),
    .Y(_07339_));
 sky130_fd_sc_hd__nand2_1 _29886_ (.A(_07322_),
    .B(_07326_),
    .Y(_07340_));
 sky130_fd_sc_hd__nor2_1 _29887_ (.A(_07339_),
    .B(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__o2bb2ai_2 _29888_ (.A1_N(_07308_),
    .A2_N(_07310_),
    .B1(_07338_),
    .B2(_07341_),
    .Y(_07342_));
 sky130_vsdinv _29889_ (.A(_07322_),
    .Y(_07343_));
 sky130_fd_sc_hd__nand2_4 _29890_ (.A(_07326_),
    .B(_07337_),
    .Y(_07344_));
 sky130_fd_sc_hd__nand2_2 _29891_ (.A(_07340_),
    .B(_07339_),
    .Y(_07345_));
 sky130_fd_sc_hd__o2111ai_4 _29892_ (.A1(_07343_),
    .A2(_07344_),
    .B1(_07345_),
    .C1(_07308_),
    .D1(_07310_),
    .Y(_07346_));
 sky130_fd_sc_hd__nand2_1 _29893_ (.A(_07342_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__nor3_4 _29894_ (.A(_06644_),
    .B(_06934_),
    .C(_07099_),
    .Y(_07348_));
 sky130_fd_sc_hd__a31oi_2 _29895_ (.A1(_07100_),
    .A2(_07133_),
    .A3(_07132_),
    .B1(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2_2 _29896_ (.A(_07347_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__nand3_1 _29897_ (.A(_07100_),
    .B(_07133_),
    .C(_07132_),
    .Y(_07351_));
 sky130_fd_sc_hd__nand2_1 _29898_ (.A(_07351_),
    .B(_07098_),
    .Y(_07352_));
 sky130_fd_sc_hd__nand3_4 _29899_ (.A(_07352_),
    .B(_07342_),
    .C(_07346_),
    .Y(_07353_));
 sky130_fd_sc_hd__buf_4 _29900_ (.A(_19872_),
    .X(_07354_));
 sky130_fd_sc_hd__nand2_1 _29901_ (.A(_07354_),
    .B(_05214_),
    .Y(_07355_));
 sky130_fd_sc_hd__buf_6 _29902_ (.A(\pcpi_mul.rs2[18] ),
    .X(_07356_));
 sky130_fd_sc_hd__nand2_2 _29903_ (.A(_07356_),
    .B(_05297_),
    .Y(_07357_));
 sky130_fd_sc_hd__nor2_2 _29904_ (.A(_07355_),
    .B(_07357_),
    .Y(_07358_));
 sky130_vsdinv _29905_ (.A(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__nand2_1 _29906_ (.A(_07355_),
    .B(_07357_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_4 _29907_ (.A(_07359_),
    .B(_07360_),
    .Y(_07361_));
 sky130_vsdinv _29908_ (.A(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__nand3_4 _29909_ (.A(_07350_),
    .B(_07353_),
    .C(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__clkbuf_4 _29910_ (.A(_07363_),
    .X(_07364_));
 sky130_fd_sc_hd__nand3_2 _29911_ (.A(_07137_),
    .B(_07142_),
    .C(_07140_),
    .Y(_07365_));
 sky130_fd_sc_hd__a21oi_2 _29912_ (.A1(_07350_),
    .A2(_07353_),
    .B1(_07362_),
    .Y(_07366_));
 sky130_fd_sc_hd__nor2_4 _29913_ (.A(_07365_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__nand2_1 _29914_ (.A(_07350_),
    .B(_07353_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand2_1 _29915_ (.A(_07368_),
    .B(_07361_),
    .Y(_07369_));
 sky130_fd_sc_hd__a21oi_4 _29916_ (.A1(_07369_),
    .A2(_07363_),
    .B1(_07144_),
    .Y(_07370_));
 sky130_fd_sc_hd__a21oi_4 _29917_ (.A1(_07364_),
    .A2(_07367_),
    .B1(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__a21oi_2 _29918_ (.A1(_07286_),
    .A2(_07288_),
    .B1(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__nor2_4 _29919_ (.A(_07150_),
    .B(_07155_),
    .Y(_07373_));
 sky130_fd_sc_hd__nand3_4 _29920_ (.A(_07286_),
    .B(_07371_),
    .C(_07288_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand3b_2 _29921_ (.A_N(_07372_),
    .B(_07373_),
    .C(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__a21oi_1 _29922_ (.A1(_07284_),
    .A2(_07280_),
    .B1(_07287_),
    .Y(_07376_));
 sky130_fd_sc_hd__nor2_1 _29923_ (.A(_07073_),
    .B(_07060_),
    .Y(_07377_));
 sky130_fd_sc_hd__o211a_1 _29924_ (.A1(_07062_),
    .A2(_07377_),
    .B1(_07280_),
    .C1(_07284_),
    .X(_07378_));
 sky130_fd_sc_hd__o21ai_2 _29925_ (.A1(_07376_),
    .A2(_07378_),
    .B1(_07371_),
    .Y(_07379_));
 sky130_fd_sc_hd__a21o_1 _29926_ (.A1(_07364_),
    .A2(_07367_),
    .B1(_07370_),
    .X(_07380_));
 sky130_fd_sc_hd__nand3_2 _29927_ (.A(_07380_),
    .B(_07286_),
    .C(_07288_),
    .Y(_07381_));
 sky130_fd_sc_hd__nand3_4 _29928_ (.A(_07379_),
    .B(_07148_),
    .C(_07381_),
    .Y(_07382_));
 sky130_vsdinv _29929_ (.A(_07013_),
    .Y(_07383_));
 sky130_fd_sc_hd__o21a_2 _29930_ (.A1(_07015_),
    .A2(_07383_),
    .B1(_07019_),
    .X(_07384_));
 sky130_fd_sc_hd__a21o_1 _29931_ (.A1(_07147_),
    .A2(_07149_),
    .B1(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__nand3_2 _29932_ (.A(_07147_),
    .B(_07149_),
    .C(_07384_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand2_1 _29933_ (.A(_07385_),
    .B(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__nand3_2 _29934_ (.A(_07375_),
    .B(_07382_),
    .C(_07387_),
    .Y(_07388_));
 sky130_vsdinv _29935_ (.A(_07145_),
    .Y(_07389_));
 sky130_fd_sc_hd__a31oi_2 _29936_ (.A1(_07075_),
    .A2(_07149_),
    .A3(_07146_),
    .B1(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand3_2 _29937_ (.A(_07374_),
    .B(_07390_),
    .C(_07077_),
    .Y(_07391_));
 sky130_fd_sc_hd__o21ai_1 _29938_ (.A1(_07372_),
    .A2(_07391_),
    .B1(_07382_),
    .Y(_07392_));
 sky130_fd_sc_hd__and2_1 _29939_ (.A(_07385_),
    .B(_07386_),
    .X(_07393_));
 sky130_fd_sc_hd__nand2_1 _29940_ (.A(_07392_),
    .B(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__o2111ai_4 _29941_ (.A1(_07161_),
    .A2(_07154_),
    .B1(_07165_),
    .C1(_07388_),
    .D1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__nand2_1 _29942_ (.A(_07153_),
    .B(_06954_),
    .Y(_07396_));
 sky130_fd_sc_hd__o22ai_4 _29943_ (.A1(_07373_),
    .A2(_07396_),
    .B1(_07161_),
    .B2(_07154_),
    .Y(_07397_));
 sky130_fd_sc_hd__nand2_1 _29944_ (.A(_07392_),
    .B(_07387_),
    .Y(_07398_));
 sky130_fd_sc_hd__nand3_2 _29945_ (.A(_07375_),
    .B(_07393_),
    .C(_07382_),
    .Y(_07399_));
 sky130_fd_sc_hd__nand3_4 _29946_ (.A(_07397_),
    .B(_07398_),
    .C(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__nand2_1 _29947_ (.A(_07395_),
    .B(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__a22oi_4 _29948_ (.A1(_07401_),
    .A2(_07159_),
    .B1(_07168_),
    .B2(_07172_),
    .Y(_07402_));
 sky130_vsdinv _29949_ (.A(_07159_),
    .Y(_07403_));
 sky130_fd_sc_hd__nand3_4 _29950_ (.A(_07395_),
    .B(_07400_),
    .C(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__and2_1 _29951_ (.A(_06894_),
    .B(_06883_),
    .X(_07405_));
 sky130_fd_sc_hd__o2bb2ai_2 _29952_ (.A1_N(_07400_),
    .A2_N(_07395_),
    .B1(_07158_),
    .B2(_07405_),
    .Y(_07406_));
 sky130_vsdinv _29953_ (.A(_07171_),
    .Y(_07407_));
 sky130_fd_sc_hd__nand2_1 _29954_ (.A(_07169_),
    .B(_07170_),
    .Y(_07408_));
 sky130_fd_sc_hd__o2bb2ai_2 _29955_ (.A1_N(_06794_),
    .A2_N(_07167_),
    .B1(_07407_),
    .B2(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__a21oi_4 _29956_ (.A1(_07406_),
    .A2(_07404_),
    .B1(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__a21oi_4 _29957_ (.A1(_07402_),
    .A2(_07404_),
    .B1(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand3_2 _29958_ (.A(_07176_),
    .B(_07177_),
    .C(_07168_),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_1 _29959_ (.A(_07184_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__xor2_1 _29960_ (.A(_07411_),
    .B(_07413_),
    .X(_02638_));
 sky130_fd_sc_hd__nor2_2 _29961_ (.A(_07372_),
    .B(_07391_),
    .Y(_07414_));
 sky130_fd_sc_hd__and3_1 _29962_ (.A(_07382_),
    .B(_07385_),
    .C(_07386_),
    .X(_07415_));
 sky130_fd_sc_hd__a22oi_4 _29963_ (.A1(_06363_),
    .A2(_05665_),
    .B1(_06895_),
    .B2(_05981_),
    .Y(_07416_));
 sky130_fd_sc_hd__buf_4 _29964_ (.A(_05294_),
    .X(_07417_));
 sky130_fd_sc_hd__and4_1 _29965_ (.A(_06363_),
    .B(_06898_),
    .C(_05696_),
    .D(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__nand2_4 _29966_ (.A(_19898_),
    .B(_05454_),
    .Y(_07419_));
 sky130_fd_sc_hd__o21ai_2 _29967_ (.A1(_07416_),
    .A2(_07418_),
    .B1(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__nand2_1 _29968_ (.A(_07102_),
    .B(_05391_),
    .Y(_07421_));
 sky130_fd_sc_hd__buf_8 _29969_ (.A(_06545_),
    .X(_07422_));
 sky130_fd_sc_hd__nand3b_4 _29970_ (.A_N(_07421_),
    .B(_07422_),
    .C(_06473_),
    .Y(_07423_));
 sky130_vsdinv _29971_ (.A(_07419_),
    .Y(_07424_));
 sky130_fd_sc_hd__a22o_1 _29972_ (.A1(_06357_),
    .A2(_06249_),
    .B1(_06607_),
    .B2(_20156_),
    .X(_07425_));
 sky130_fd_sc_hd__nand3_2 _29973_ (.A(_07423_),
    .B(_07424_),
    .C(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__o21ai_2 _29974_ (.A1(_07316_),
    .A2(_07312_),
    .B1(_07318_),
    .Y(_07427_));
 sky130_fd_sc_hd__nand3_4 _29975_ (.A(_07420_),
    .B(_07426_),
    .C(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__o21ai_2 _29976_ (.A1(_07416_),
    .A2(_07418_),
    .B1(_07424_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand3_2 _29977_ (.A(_07423_),
    .B(_07419_),
    .C(_07425_),
    .Y(_07430_));
 sky130_fd_sc_hd__a21oi_2 _29978_ (.A1(_07319_),
    .A2(_07320_),
    .B1(_07315_),
    .Y(_07431_));
 sky130_fd_sc_hd__nand3_4 _29979_ (.A(_07429_),
    .B(_07430_),
    .C(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__a22oi_4 _29980_ (.A1(_06118_),
    .A2(_06289_),
    .B1(_06045_),
    .B2(_20146_),
    .Y(_07433_));
 sky130_fd_sc_hd__nand2_2 _29981_ (.A(_06041_),
    .B(_05689_),
    .Y(_07434_));
 sky130_fd_sc_hd__nand2_2 _29982_ (.A(_06534_),
    .B(_07033_),
    .Y(_07435_));
 sky130_fd_sc_hd__nor2_4 _29983_ (.A(_07434_),
    .B(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__nand2_2 _29984_ (.A(_19909_),
    .B(_20142_),
    .Y(_07437_));
 sky130_fd_sc_hd__o21bai_2 _29985_ (.A1(_07433_),
    .A2(_07436_),
    .B1_N(_07437_),
    .Y(_07438_));
 sky130_fd_sc_hd__nand3b_4 _29986_ (.A_N(_07434_),
    .B(_07333_),
    .C(_05823_),
    .Y(_07439_));
 sky130_fd_sc_hd__nand2_2 _29987_ (.A(_07434_),
    .B(_07435_),
    .Y(_07440_));
 sky130_fd_sc_hd__nand3_2 _29988_ (.A(_07439_),
    .B(_07437_),
    .C(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__nand2_4 _29989_ (.A(_07438_),
    .B(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__nand3_1 _29990_ (.A(_07428_),
    .B(_07432_),
    .C(_07442_),
    .Y(_07443_));
 sky130_vsdinv _29991_ (.A(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__a21oi_4 _29992_ (.A1(_07428_),
    .A2(_07432_),
    .B1(_07442_),
    .Y(_07445_));
 sky130_fd_sc_hd__buf_4 _29993_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07446_));
 sky130_fd_sc_hd__nand3_4 _29994_ (.A(_07446_),
    .B(_19886_),
    .C(_05176_),
    .Y(_07447_));
 sky130_fd_sc_hd__nor2_8 _29995_ (.A(_05252_),
    .B(_07447_),
    .Y(_07448_));
 sky130_fd_sc_hd__buf_6 _29996_ (.A(_07089_),
    .X(_07449_));
 sky130_fd_sc_hd__a22o_2 _29997_ (.A1(_07088_),
    .A2(_05245_),
    .B1(_07449_),
    .B2(_06199_),
    .X(_07450_));
 sky130_fd_sc_hd__nand2_4 _29998_ (.A(_06640_),
    .B(_20162_),
    .Y(_07451_));
 sky130_vsdinv _29999_ (.A(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand2_1 _30000_ (.A(_07450_),
    .B(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__a22oi_4 _30001_ (.A1(_07289_),
    .A2(_05245_),
    .B1(_07449_),
    .B2(_05244_),
    .Y(_07454_));
 sky130_fd_sc_hd__o21ai_2 _30002_ (.A1(_07454_),
    .A2(_07448_),
    .B1(_07451_),
    .Y(_07455_));
 sky130_fd_sc_hd__o211ai_4 _30003_ (.A1(_07448_),
    .A2(_07453_),
    .B1(_07358_),
    .C1(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__o21ai_2 _30004_ (.A1(_07454_),
    .A2(_07448_),
    .B1(_07452_),
    .Y(_07457_));
 sky130_fd_sc_hd__o211ai_4 _30005_ (.A1(_05253_),
    .A2(_07447_),
    .B1(_07451_),
    .C1(_07450_),
    .Y(_07458_));
 sky130_fd_sc_hd__nand3_4 _30006_ (.A(_07457_),
    .B(_07359_),
    .C(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__nor2_2 _30007_ (.A(_07302_),
    .B(_07301_),
    .Y(_07460_));
 sky130_fd_sc_hd__nor2_4 _30008_ (.A(_07296_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__a21o_2 _30009_ (.A1(_07456_),
    .A2(_07459_),
    .B1(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__nand3_4 _30010_ (.A(_07456_),
    .B(_07459_),
    .C(_07461_),
    .Y(_07463_));
 sky130_vsdinv _30011_ (.A(_07307_),
    .Y(_07464_));
 sky130_fd_sc_hd__a21oi_4 _30012_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__nand2_2 _30013_ (.A(_07459_),
    .B(_07461_),
    .Y(_07466_));
 sky130_vsdinv _30014_ (.A(_07456_),
    .Y(_07467_));
 sky130_fd_sc_hd__o211a_1 _30015_ (.A1(_07466_),
    .A2(_07467_),
    .B1(_07464_),
    .C1(_07462_),
    .X(_07468_));
 sky130_fd_sc_hd__o22ai_4 _30016_ (.A1(_07444_),
    .A2(_07445_),
    .B1(_07465_),
    .B2(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__a21o_1 _30017_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07464_),
    .X(_07470_));
 sky130_fd_sc_hd__nand3_4 _30018_ (.A(_07462_),
    .B(_07464_),
    .C(_07463_),
    .Y(_07471_));
 sky130_fd_sc_hd__nor2_4 _30019_ (.A(_07445_),
    .B(_07444_),
    .Y(_07472_));
 sky130_fd_sc_hd__nand3_4 _30020_ (.A(_07470_),
    .B(_07471_),
    .C(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__nand2_4 _30021_ (.A(_07346_),
    .B(_07308_),
    .Y(_07474_));
 sky130_fd_sc_hd__a21oi_4 _30022_ (.A1(_07469_),
    .A2(_07473_),
    .B1(_07474_),
    .Y(_07475_));
 sky130_vsdinv _30023_ (.A(_07308_),
    .Y(_07476_));
 sky130_fd_sc_hd__o2111a_1 _30024_ (.A1(_07343_),
    .A2(_07344_),
    .B1(_07345_),
    .C1(_07308_),
    .D1(_07310_),
    .X(_07477_));
 sky130_fd_sc_hd__o211a_2 _30025_ (.A1(_07476_),
    .A2(_07477_),
    .B1(_07473_),
    .C1(_07469_),
    .X(_07478_));
 sky130_fd_sc_hd__buf_8 _30026_ (.A(_07356_),
    .X(_07479_));
 sky130_fd_sc_hd__nand2_4 _30027_ (.A(_07479_),
    .B(_05144_),
    .Y(_07480_));
 sky130_fd_sc_hd__buf_4 _30028_ (.A(\pcpi_mul.rs2[20] ),
    .X(_07481_));
 sky130_fd_sc_hd__buf_6 _30029_ (.A(_07481_),
    .X(_07482_));
 sky130_fd_sc_hd__buf_6 _30030_ (.A(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__a22oi_4 _30031_ (.A1(_07483_),
    .A2(_05415_),
    .B1(_19874_),
    .B2(_05147_),
    .Y(_07484_));
 sky130_fd_sc_hd__nand2_2 _30032_ (.A(_07354_),
    .B(_05297_),
    .Y(_07485_));
 sky130_fd_sc_hd__nand2_2 _30033_ (.A(_07482_),
    .B(_05214_),
    .Y(_07486_));
 sky130_fd_sc_hd__nor2_4 _30034_ (.A(_07485_),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__nor2_4 _30035_ (.A(_07484_),
    .B(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__xor2_4 _30036_ (.A(_07480_),
    .B(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__o21ai_4 _30037_ (.A1(_07475_),
    .A2(_07478_),
    .B1(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__nand2_2 _30038_ (.A(_07469_),
    .B(_07473_),
    .Y(_07491_));
 sky130_vsdinv _30039_ (.A(_07474_),
    .Y(_07492_));
 sky130_fd_sc_hd__nand2_2 _30040_ (.A(_07491_),
    .B(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__nand3_4 _30041_ (.A(_07469_),
    .B(_07474_),
    .C(_07473_),
    .Y(_07494_));
 sky130_fd_sc_hd__nand3b_4 _30042_ (.A_N(_07489_),
    .B(_07493_),
    .C(_07494_),
    .Y(_07495_));
 sky130_vsdinv _30043_ (.A(_07364_),
    .Y(_07496_));
 sky130_fd_sc_hd__a21oi_4 _30044_ (.A1(_07490_),
    .A2(_07495_),
    .B1(_07496_),
    .Y(_07497_));
 sky130_fd_sc_hd__nand3_4 _30045_ (.A(_07490_),
    .B(_07496_),
    .C(_07495_),
    .Y(_07498_));
 sky130_vsdinv _30046_ (.A(_07498_),
    .Y(_07499_));
 sky130_vsdinv _30047_ (.A(_07200_),
    .Y(_07500_));
 sky130_fd_sc_hd__nor2_2 _30048_ (.A(_07203_),
    .B(_07209_),
    .Y(_07501_));
 sky130_fd_sc_hd__buf_6 _30049_ (.A(_20137_),
    .X(_07502_));
 sky130_fd_sc_hd__buf_6 _30050_ (.A(_06441_),
    .X(_07503_));
 sky130_fd_sc_hd__a22oi_4 _30051_ (.A1(_06478_),
    .A2(_07502_),
    .B1(_06097_),
    .B2(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand3_4 _30052_ (.A(_19911_),
    .B(_06110_),
    .C(_06309_),
    .Y(_07505_));
 sky130_fd_sc_hd__nor2_8 _30053_ (.A(_06722_),
    .B(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_2 _30054_ (.A(_19917_),
    .B(_06989_),
    .Y(_07507_));
 sky130_fd_sc_hd__o21ai_2 _30055_ (.A1(_07504_),
    .A2(_07506_),
    .B1(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__o21ai_2 _30056_ (.A1(_07331_),
    .A2(_07327_),
    .B1(_07334_),
    .Y(_07509_));
 sky130_fd_sc_hd__buf_8 _30057_ (.A(_06722_),
    .X(_07510_));
 sky130_vsdinv _30058_ (.A(_07507_),
    .Y(_07511_));
 sky130_fd_sc_hd__a22o_2 _30059_ (.A1(_06095_),
    .A2(_20138_),
    .B1(_06657_),
    .B2(_07503_),
    .X(_07512_));
 sky130_fd_sc_hd__o211ai_4 _30060_ (.A1(_07510_),
    .A2(_07505_),
    .B1(_07511_),
    .C1(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand3_4 _30061_ (.A(_07508_),
    .B(_07509_),
    .C(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__o21ai_2 _30062_ (.A1(_07504_),
    .A2(_07506_),
    .B1(_07511_),
    .Y(_07515_));
 sky130_vsdinv _30063_ (.A(_07331_),
    .Y(_07516_));
 sky130_fd_sc_hd__a21oi_2 _30064_ (.A1(_07516_),
    .A2(_07335_),
    .B1(_07330_),
    .Y(_07517_));
 sky130_fd_sc_hd__o211ai_4 _30065_ (.A1(_07510_),
    .A2(_07505_),
    .B1(_07507_),
    .C1(_07512_),
    .Y(_07518_));
 sky130_fd_sc_hd__nand3_4 _30066_ (.A(_07515_),
    .B(_07517_),
    .C(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__nor2_8 _30067_ (.A(_07192_),
    .B(_07188_),
    .Y(_07520_));
 sky130_fd_sc_hd__o2bb2ai_4 _30068_ (.A1_N(_07514_),
    .A2_N(_07519_),
    .B1(_07186_),
    .B2(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__nor2_4 _30069_ (.A(_07186_),
    .B(_07520_),
    .Y(_07522_));
 sky130_fd_sc_hd__nand3_4 _30070_ (.A(_07519_),
    .B(_07514_),
    .C(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__nand2_4 _30071_ (.A(_07344_),
    .B(_07322_),
    .Y(_07524_));
 sky130_fd_sc_hd__a21oi_4 _30072_ (.A1(_07521_),
    .A2(_07523_),
    .B1(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__nand2_1 _30073_ (.A(_07519_),
    .B(_07522_),
    .Y(_07526_));
 sky130_vsdinv _30074_ (.A(_07514_),
    .Y(_07527_));
 sky130_fd_sc_hd__o211a_1 _30075_ (.A1(_07526_),
    .A2(_07527_),
    .B1(_07521_),
    .C1(_07524_),
    .X(_07528_));
 sky130_fd_sc_hd__o22ai_4 _30076_ (.A1(_07500_),
    .A2(_07501_),
    .B1(_07525_),
    .B2(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__and2_1 _30077_ (.A(_07208_),
    .B(_07196_),
    .X(_07530_));
 sky130_fd_sc_hd__nand2_1 _30078_ (.A(_07521_),
    .B(_07523_),
    .Y(_07531_));
 sky130_fd_sc_hd__and2_1 _30079_ (.A(_07344_),
    .B(_07322_),
    .X(_07532_));
 sky130_fd_sc_hd__nand2_2 _30080_ (.A(_07531_),
    .B(_07532_),
    .Y(_07533_));
 sky130_fd_sc_hd__nand3_4 _30081_ (.A(_07524_),
    .B(_07521_),
    .C(_07523_),
    .Y(_07534_));
 sky130_fd_sc_hd__nand3b_4 _30082_ (.A_N(_07530_),
    .B(_07533_),
    .C(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__o21ai_4 _30083_ (.A1(_07222_),
    .A2(_07207_),
    .B1(_07216_),
    .Y(_07536_));
 sky130_fd_sc_hd__a21oi_4 _30084_ (.A1(_07529_),
    .A2(_07535_),
    .B1(_07536_),
    .Y(_07537_));
 sky130_vsdinv _30085_ (.A(_07204_),
    .Y(_07538_));
 sky130_fd_sc_hd__o2bb2ai_1 _30086_ (.A1_N(_07532_),
    .A2_N(_07531_),
    .B1(_07209_),
    .B2(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__o211a_2 _30087_ (.A1(_07528_),
    .A2(_07539_),
    .B1(_07536_),
    .C1(_07529_),
    .X(_07540_));
 sky130_fd_sc_hd__nor2_8 _30088_ (.A(_07252_),
    .B(_07255_),
    .Y(_07541_));
 sky130_fd_sc_hd__a21boi_2 _30089_ (.A1(_07262_),
    .A2(_07247_),
    .B1_N(_07243_),
    .Y(_07542_));
 sky130_fd_sc_hd__buf_6 _30090_ (.A(_06701_),
    .X(_07543_));
 sky130_fd_sc_hd__a22oi_4 _30091_ (.A1(_19920_),
    .A2(_06714_),
    .B1(_05674_),
    .B2(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__nand2_4 _30092_ (.A(_06986_),
    .B(net473),
    .Y(_07545_));
 sky130_fd_sc_hd__nand2_4 _30093_ (.A(_05377_),
    .B(_07257_),
    .Y(_07546_));
 sky130_fd_sc_hd__nor2_8 _30094_ (.A(_07545_),
    .B(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__buf_6 _30095_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07548_));
 sky130_fd_sc_hd__nand2_4 _30096_ (.A(net469),
    .B(_07548_),
    .Y(_07549_));
 sky130_vsdinv _30097_ (.A(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__o21ai_2 _30098_ (.A1(_07544_),
    .A2(_07547_),
    .B1(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__or2_2 _30099_ (.A(_07545_),
    .B(_07546_),
    .X(_07552_));
 sky130_fd_sc_hd__nand2_4 _30100_ (.A(_07545_),
    .B(_07546_),
    .Y(_07553_));
 sky130_fd_sc_hd__nand3_2 _30101_ (.A(_07552_),
    .B(_07553_),
    .C(_07549_),
    .Y(_07554_));
 sky130_fd_sc_hd__o2111ai_4 _30102_ (.A1(_07235_),
    .A2(_07234_),
    .B1(_07239_),
    .C1(_07551_),
    .D1(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__nand3_4 _30103_ (.A(_07552_),
    .B(_07553_),
    .C(_07550_),
    .Y(_07556_));
 sky130_fd_sc_hd__o21ai_4 _30104_ (.A1(_07235_),
    .A2(_07234_),
    .B1(_07239_),
    .Y(_07557_));
 sky130_fd_sc_hd__o21ai_4 _30105_ (.A1(_07544_),
    .A2(_07547_),
    .B1(_07549_),
    .Y(_07558_));
 sky130_fd_sc_hd__nand3_4 _30106_ (.A(_07556_),
    .B(_07557_),
    .C(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand2_1 _30107_ (.A(_07555_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__buf_6 _30108_ (.A(_20113_),
    .X(_07561_));
 sky130_fd_sc_hd__nand2_1 _30109_ (.A(_19931_),
    .B(_20118_),
    .Y(_07562_));
 sky130_fd_sc_hd__a21o_1 _30110_ (.A1(_05821_),
    .A2(_07561_),
    .B1(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__buf_4 _30111_ (.A(_07232_),
    .X(_07564_));
 sky130_fd_sc_hd__nand2_1 _30112_ (.A(_05284_),
    .B(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__a21o_1 _30113_ (.A1(_05236_),
    .A2(_07250_),
    .B1(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__buf_4 _30114_ (.A(_20122_),
    .X(_07567_));
 sky130_fd_sc_hd__buf_4 _30115_ (.A(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__nand2_2 _30116_ (.A(_05830_),
    .B(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__a21o_4 _30117_ (.A1(_07563_),
    .A2(_07566_),
    .B1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__nand3_4 _30118_ (.A(_07563_),
    .B(_07566_),
    .C(_07569_),
    .Y(_07571_));
 sky130_fd_sc_hd__and2_1 _30119_ (.A(_07570_),
    .B(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__nand2_1 _30120_ (.A(_07560_),
    .B(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__nand2_2 _30121_ (.A(_07570_),
    .B(_07571_),
    .Y(_07574_));
 sky130_fd_sc_hd__nand3_2 _30122_ (.A(_07555_),
    .B(_07574_),
    .C(_07559_),
    .Y(_07575_));
 sky130_fd_sc_hd__nand3_4 _30123_ (.A(_07542_),
    .B(_07573_),
    .C(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__o21a_1 _30124_ (.A1(_07541_),
    .A2(_07260_),
    .B1(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__a21bo_1 _30125_ (.A1(_07262_),
    .A2(_07247_),
    .B1_N(_07243_),
    .X(_07578_));
 sky130_fd_sc_hd__nand3_2 _30126_ (.A(_07572_),
    .B(_07555_),
    .C(_07559_),
    .Y(_07579_));
 sky130_fd_sc_hd__nand2_1 _30127_ (.A(_07560_),
    .B(_07574_),
    .Y(_07580_));
 sky130_fd_sc_hd__nand3_4 _30128_ (.A(_07578_),
    .B(_07579_),
    .C(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__nor2_1 _30129_ (.A(_07541_),
    .B(_07260_),
    .Y(_07582_));
 sky130_vsdinv _30130_ (.A(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__a21oi_4 _30131_ (.A1(_07581_),
    .A2(_07576_),
    .B1(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__a21oi_4 _30132_ (.A1(_07577_),
    .A2(_07581_),
    .B1(_07584_),
    .Y(_07585_));
 sky130_fd_sc_hd__o21ai_2 _30133_ (.A1(_07537_),
    .A2(_07540_),
    .B1(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__a21o_1 _30134_ (.A1(_07529_),
    .A2(_07535_),
    .B1(_07536_),
    .X(_07587_));
 sky130_fd_sc_hd__a21o_1 _30135_ (.A1(_07581_),
    .A2(_07576_),
    .B1(_07583_),
    .X(_07588_));
 sky130_fd_sc_hd__nand3_1 _30136_ (.A(_07581_),
    .B(_07576_),
    .C(_07583_),
    .Y(_07589_));
 sky130_fd_sc_hd__nand2_1 _30137_ (.A(_07588_),
    .B(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__nand3_4 _30138_ (.A(_07529_),
    .B(_07535_),
    .C(_07536_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand3_2 _30139_ (.A(_07587_),
    .B(_07590_),
    .C(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__nand3_4 _30140_ (.A(_07586_),
    .B(_07353_),
    .C(_07592_),
    .Y(_07593_));
 sky130_vsdinv _30141_ (.A(_07589_),
    .Y(_07594_));
 sky130_fd_sc_hd__o22ai_4 _30142_ (.A1(_07594_),
    .A2(_07584_),
    .B1(_07537_),
    .B2(_07540_),
    .Y(_07595_));
 sky130_vsdinv _30143_ (.A(_07353_),
    .Y(_07596_));
 sky130_fd_sc_hd__nand3_4 _30144_ (.A(_07587_),
    .B(_07585_),
    .C(_07591_),
    .Y(_07597_));
 sky130_fd_sc_hd__nand3_4 _30145_ (.A(_07595_),
    .B(_07596_),
    .C(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__a21bo_2 _30146_ (.A1(_07278_),
    .A2(_07224_),
    .B1_N(_07218_),
    .X(_07599_));
 sky130_fd_sc_hd__a21oi_4 _30147_ (.A1(_07593_),
    .A2(_07598_),
    .B1(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__and3_1 _30148_ (.A(_07593_),
    .B(_07598_),
    .C(_07599_),
    .X(_07601_));
 sky130_fd_sc_hd__o22ai_4 _30149_ (.A1(_07497_),
    .A2(_07499_),
    .B1(_07600_),
    .B2(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__nand2_2 _30150_ (.A(_07493_),
    .B(_07494_),
    .Y(_07603_));
 sky130_fd_sc_hd__a21oi_1 _30151_ (.A1(_07603_),
    .A2(_07489_),
    .B1(_07364_),
    .Y(_07604_));
 sky130_fd_sc_hd__a21oi_2 _30152_ (.A1(_07495_),
    .A2(_07604_),
    .B1(_07497_),
    .Y(_07605_));
 sky130_fd_sc_hd__a21o_1 _30153_ (.A1(_07593_),
    .A2(_07598_),
    .B1(_07599_),
    .X(_07606_));
 sky130_fd_sc_hd__nand3_4 _30154_ (.A(_07593_),
    .B(_07598_),
    .C(_07599_),
    .Y(_07607_));
 sky130_fd_sc_hd__nand3_4 _30155_ (.A(_07605_),
    .B(_07606_),
    .C(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__nand2_1 _30156_ (.A(_07367_),
    .B(_07364_),
    .Y(_07609_));
 sky130_fd_sc_hd__nand2_4 _30157_ (.A(_07374_),
    .B(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__a21o_1 _30158_ (.A1(_07602_),
    .A2(_07608_),
    .B1(_07610_),
    .X(_07611_));
 sky130_fd_sc_hd__nor2b_4 _30159_ (.A(_07277_),
    .B_N(_07271_),
    .Y(_07612_));
 sky130_fd_sc_hd__and3_1 _30160_ (.A(_07288_),
    .B(_07280_),
    .C(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__nand2_2 _30161_ (.A(_07288_),
    .B(_07280_),
    .Y(_07614_));
 sky130_vsdinv _30162_ (.A(_07614_),
    .Y(_07615_));
 sky130_fd_sc_hd__nor2_8 _30163_ (.A(_07612_),
    .B(_07615_),
    .Y(_07616_));
 sky130_fd_sc_hd__nor2_2 _30164_ (.A(_07613_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__nand3_4 _30165_ (.A(_07602_),
    .B(_07610_),
    .C(_07608_),
    .Y(_07618_));
 sky130_fd_sc_hd__nand3_4 _30166_ (.A(_07611_),
    .B(_07617_),
    .C(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__a21oi_4 _30167_ (.A1(_07602_),
    .A2(_07608_),
    .B1(_07610_),
    .Y(_07620_));
 sky130_fd_sc_hd__o2bb2ai_2 _30168_ (.A1_N(_07490_),
    .A2_N(_07495_),
    .B1(_07368_),
    .B2(_07361_),
    .Y(_07621_));
 sky130_fd_sc_hd__nand3_4 _30169_ (.A(_07607_),
    .B(_07621_),
    .C(_07498_),
    .Y(_07622_));
 sky130_fd_sc_hd__o211a_1 _30170_ (.A1(_07600_),
    .A2(_07622_),
    .B1(_07610_),
    .C1(_07602_),
    .X(_07623_));
 sky130_fd_sc_hd__o22ai_4 _30171_ (.A1(_07616_),
    .A2(_07613_),
    .B1(_07620_),
    .B2(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__o211a_2 _30172_ (.A1(_07414_),
    .A2(_07415_),
    .B1(_07619_),
    .C1(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__nand2_1 _30173_ (.A(_07624_),
    .B(_07619_),
    .Y(_07626_));
 sky130_fd_sc_hd__nor2_1 _30174_ (.A(_07414_),
    .B(_07415_),
    .Y(_07627_));
 sky130_fd_sc_hd__nand2_2 _30175_ (.A(_07626_),
    .B(_07627_),
    .Y(_07628_));
 sky130_vsdinv _30176_ (.A(_07385_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand2_4 _30177_ (.A(_07628_),
    .B(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__nor2_1 _30178_ (.A(_07625_),
    .B(_07630_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_1 _30179_ (.A(_07147_),
    .B(_07149_),
    .Y(_07632_));
 sky130_vsdinv _30180_ (.A(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__a21o_1 _30181_ (.A1(_07393_),
    .A2(_07382_),
    .B1(_07414_),
    .X(_07634_));
 sky130_fd_sc_hd__a21oi_4 _30182_ (.A1(_07624_),
    .A2(_07619_),
    .B1(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__o22ai_4 _30183_ (.A1(_07384_),
    .A2(_07633_),
    .B1(_07635_),
    .B2(_07625_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand2_1 _30184_ (.A(_07395_),
    .B(_07403_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_2 _30185_ (.A(_07637_),
    .B(_07400_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _30186_ (.A(_07636_),
    .B(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__o21ai_1 _30187_ (.A1(_07635_),
    .A2(_07625_),
    .B1(_07629_),
    .Y(_07640_));
 sky130_fd_sc_hd__nand3_4 _30188_ (.A(_07624_),
    .B(_07634_),
    .C(_07619_),
    .Y(_07641_));
 sky130_fd_sc_hd__nand3_1 _30189_ (.A(_07628_),
    .B(_07385_),
    .C(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__nand3b_2 _30190_ (.A_N(_07638_),
    .B(_07640_),
    .C(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__o21a_2 _30191_ (.A1(_07631_),
    .A2(_07639_),
    .B1(_07643_),
    .X(_07644_));
 sky130_vsdinv _30192_ (.A(_06969_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand2_2 _30193_ (.A(_06967_),
    .B(_06968_),
    .Y(_07646_));
 sky130_fd_sc_hd__a21oi_2 _30194_ (.A1(_07645_),
    .A2(_07646_),
    .B1(_06788_),
    .Y(_07647_));
 sky130_fd_sc_hd__o2111ai_4 _30195_ (.A1(_07645_),
    .A2(_07646_),
    .B1(_07411_),
    .C1(_07647_),
    .D1(_07179_),
    .Y(_07648_));
 sky130_fd_sc_hd__or2b_1 _30196_ (.A(_07648_),
    .B_N(_06601_),
    .X(_07649_));
 sky130_fd_sc_hd__o2bb2ai_2 _30197_ (.A1_N(_07404_),
    .A2_N(_07402_),
    .B1(_07412_),
    .B2(_07410_),
    .Y(_07650_));
 sky130_fd_sc_hd__a31oi_4 _30198_ (.A1(_07179_),
    .A2(_07181_),
    .A3(_07411_),
    .B1(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__and2_1 _30199_ (.A(_07649_),
    .B(_07651_),
    .X(_07652_));
 sky130_fd_sc_hd__xnor2_2 _30200_ (.A(_07644_),
    .B(_07652_),
    .Y(_02639_));
 sky130_fd_sc_hd__o211ai_4 _30201_ (.A1(_07625_),
    .A2(_07630_),
    .B1(_07638_),
    .C1(_07636_),
    .Y(_07653_));
 sky130_fd_sc_hd__nand2_1 _30202_ (.A(_07652_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__xor2_4 _30203_ (.A(_07612_),
    .B(_07614_),
    .X(_07655_));
 sky130_fd_sc_hd__nand2_1 _30204_ (.A(_07490_),
    .B(_07495_),
    .Y(_07656_));
 sky130_fd_sc_hd__o22ai_4 _30205_ (.A1(_07364_),
    .A2(_07656_),
    .B1(_07600_),
    .B2(_07622_),
    .Y(_07657_));
 sky130_fd_sc_hd__and2_2 _30206_ (.A(_07519_),
    .B(_07522_),
    .X(_07658_));
 sky130_fd_sc_hd__a22oi_4 _30207_ (.A1(_06100_),
    .A2(_06143_),
    .B1(_06474_),
    .B2(_06718_),
    .Y(_07659_));
 sky130_fd_sc_hd__buf_6 _30208_ (.A(\pcpi_mul.rs2[8] ),
    .X(_07660_));
 sky130_fd_sc_hd__buf_8 _30209_ (.A(\pcpi_mul.rs1[13] ),
    .X(_07661_));
 sky130_fd_sc_hd__nand3_4 _30210_ (.A(_07660_),
    .B(_06840_),
    .C(_07661_),
    .Y(_07662_));
 sky130_fd_sc_hd__nor2_2 _30211_ (.A(_06440_),
    .B(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__nand2_2 _30212_ (.A(_19917_),
    .B(_06813_),
    .Y(_07664_));
 sky130_fd_sc_hd__o21ai_2 _30213_ (.A1(_07659_),
    .A2(_07663_),
    .B1(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__o21ai_2 _30214_ (.A1(_07437_),
    .A2(_07433_),
    .B1(_07439_),
    .Y(_07666_));
 sky130_vsdinv _30215_ (.A(_07664_),
    .Y(_07667_));
 sky130_fd_sc_hd__a22o_2 _30216_ (.A1(_06483_),
    .A2(_20135_),
    .B1(_06474_),
    .B2(_20133_),
    .X(_07668_));
 sky130_fd_sc_hd__o211ai_4 _30217_ (.A1(_06452_),
    .A2(_07662_),
    .B1(_07667_),
    .C1(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__nand3_4 _30218_ (.A(_07665_),
    .B(_07666_),
    .C(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__a31oi_4 _30219_ (.A1(_07440_),
    .A2(_19910_),
    .A3(_20143_),
    .B1(_07436_),
    .Y(_07671_));
 sky130_fd_sc_hd__o21ai_2 _30220_ (.A1(_07659_),
    .A2(_07663_),
    .B1(_07667_),
    .Y(_07672_));
 sky130_fd_sc_hd__o211ai_2 _30221_ (.A1(_06452_),
    .A2(_07662_),
    .B1(_07664_),
    .C1(_07668_),
    .Y(_07673_));
 sky130_fd_sc_hd__nand3_4 _30222_ (.A(_07671_),
    .B(_07672_),
    .C(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__nor2_8 _30223_ (.A(_07511_),
    .B(_07506_),
    .Y(_07675_));
 sky130_fd_sc_hd__o2bb2ai_4 _30224_ (.A1_N(_07670_),
    .A2_N(_07674_),
    .B1(_07504_),
    .B2(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__nor2_4 _30225_ (.A(_07504_),
    .B(_07675_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand3_4 _30226_ (.A(_07674_),
    .B(_07670_),
    .C(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand2_1 _30227_ (.A(_07432_),
    .B(_07442_),
    .Y(_07679_));
 sky130_fd_sc_hd__nand2_4 _30228_ (.A(_07679_),
    .B(_07428_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21oi_4 _30229_ (.A1(_07676_),
    .A2(_07678_),
    .B1(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__and3_1 _30230_ (.A(_07665_),
    .B(_07666_),
    .C(_07669_),
    .X(_07682_));
 sky130_fd_sc_hd__nand2_1 _30231_ (.A(_07674_),
    .B(_07677_),
    .Y(_07683_));
 sky130_fd_sc_hd__o211a_2 _30232_ (.A1(_07682_),
    .A2(_07683_),
    .B1(_07676_),
    .C1(_07680_),
    .X(_07684_));
 sky130_fd_sc_hd__o22ai_4 _30233_ (.A1(_07527_),
    .A2(_07658_),
    .B1(_07681_),
    .B2(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__nand2_1 _30234_ (.A(_07534_),
    .B(_07530_),
    .Y(_07686_));
 sky130_fd_sc_hd__nand2_1 _30235_ (.A(_07686_),
    .B(_07533_),
    .Y(_07687_));
 sky130_fd_sc_hd__a21o_1 _30236_ (.A1(_07676_),
    .A2(_07678_),
    .B1(_07680_),
    .X(_07688_));
 sky130_fd_sc_hd__nand3_4 _30237_ (.A(_07680_),
    .B(_07676_),
    .C(_07678_),
    .Y(_07689_));
 sky130_fd_sc_hd__nor2_4 _30238_ (.A(_07527_),
    .B(_07658_),
    .Y(_07690_));
 sky130_fd_sc_hd__nand3_2 _30239_ (.A(_07688_),
    .B(_07689_),
    .C(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__nand3_4 _30240_ (.A(_07685_),
    .B(_07687_),
    .C(_07691_),
    .Y(_07692_));
 sky130_vsdinv _30241_ (.A(_07519_),
    .Y(_07693_));
 sky130_fd_sc_hd__nor2_2 _30242_ (.A(_07522_),
    .B(_07527_),
    .Y(_07694_));
 sky130_fd_sc_hd__o22ai_4 _30243_ (.A1(_07693_),
    .A2(_07694_),
    .B1(_07681_),
    .B2(_07684_),
    .Y(_07695_));
 sky130_fd_sc_hd__o21ai_2 _30244_ (.A1(_07530_),
    .A2(_07525_),
    .B1(_07534_),
    .Y(_07696_));
 sky130_fd_sc_hd__o211ai_2 _30245_ (.A1(_07527_),
    .A2(_07658_),
    .B1(_07689_),
    .C1(_07688_),
    .Y(_07697_));
 sky130_fd_sc_hd__nand3_4 _30246_ (.A(_07695_),
    .B(_07696_),
    .C(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand2_1 _30247_ (.A(_07692_),
    .B(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__or2_4 _30248_ (.A(_07562_),
    .B(_07565_),
    .X(_07700_));
 sky130_fd_sc_hd__nand2_2 _30249_ (.A(_06986_),
    .B(_07257_),
    .Y(_07701_));
 sky130_fd_sc_hd__buf_4 _30250_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07702_));
 sky130_fd_sc_hd__nand2_2 _30251_ (.A(_05377_),
    .B(_07702_),
    .Y(_07703_));
 sky130_fd_sc_hd__or2_2 _30252_ (.A(_07701_),
    .B(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__nand2_1 _30253_ (.A(_07701_),
    .B(_07703_),
    .Y(_07705_));
 sky130_fd_sc_hd__nand2_4 _30254_ (.A(_05192_),
    .B(_20107_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand3_2 _30255_ (.A(_07704_),
    .B(_07705_),
    .C(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__a21oi_4 _30256_ (.A1(_07550_),
    .A2(_07553_),
    .B1(_07547_),
    .Y(_07708_));
 sky130_fd_sc_hd__buf_4 _30257_ (.A(\pcpi_mul.rs1[16] ),
    .X(_07709_));
 sky130_fd_sc_hd__a22oi_4 _30258_ (.A1(_05797_),
    .A2(_07709_),
    .B1(_19925_),
    .B2(_07567_),
    .Y(_07710_));
 sky130_fd_sc_hd__nor2_4 _30259_ (.A(_07701_),
    .B(_07703_),
    .Y(_07711_));
 sky130_fd_sc_hd__o21bai_2 _30260_ (.A1(_07710_),
    .A2(_07711_),
    .B1_N(_07706_),
    .Y(_07712_));
 sky130_fd_sc_hd__nand3_4 _30261_ (.A(_07707_),
    .B(_07708_),
    .C(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__nor2_1 _30262_ (.A(_07706_),
    .B(_07710_),
    .Y(_07714_));
 sky130_fd_sc_hd__nand2_1 _30263_ (.A(_07714_),
    .B(_07704_),
    .Y(_07715_));
 sky130_fd_sc_hd__o21ai_2 _30264_ (.A1(_07710_),
    .A2(_07711_),
    .B1(_07706_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand3b_4 _30265_ (.A_N(_07708_),
    .B(_07715_),
    .C(_07716_),
    .Y(_07717_));
 sky130_vsdinv _30266_ (.A(_07254_),
    .Y(_07718_));
 sky130_fd_sc_hd__nand2_2 _30267_ (.A(_05141_),
    .B(_07548_),
    .Y(_07719_));
 sky130_fd_sc_hd__nand3_4 _30268_ (.A(_07719_),
    .B(_06314_),
    .C(_07561_),
    .Y(_07720_));
 sky130_fd_sc_hd__nand2_2 _30269_ (.A(_05139_),
    .B(_07233_),
    .Y(_07721_));
 sky130_fd_sc_hd__clkbuf_4 _30270_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07722_));
 sky130_fd_sc_hd__clkbuf_8 _30271_ (.A(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__nand3_4 _30272_ (.A(_07721_),
    .B(_05821_),
    .C(_07723_),
    .Y(_07724_));
 sky130_fd_sc_hd__o211a_2 _30273_ (.A1(_05186_),
    .A2(_07718_),
    .B1(_07720_),
    .C1(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__buf_4 _30274_ (.A(_07254_),
    .X(_07726_));
 sky130_fd_sc_hd__nand2_1 _30275_ (.A(_05830_),
    .B(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__a21oi_4 _30276_ (.A1(_07720_),
    .A2(_07724_),
    .B1(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__o2bb2ai_4 _30277_ (.A1_N(_07713_),
    .A2_N(_07717_),
    .B1(_07725_),
    .B2(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__nor2_2 _30278_ (.A(_07728_),
    .B(_07725_),
    .Y(_07730_));
 sky130_fd_sc_hd__nand3_4 _30279_ (.A(_07717_),
    .B(_07713_),
    .C(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__a21oi_4 _30280_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_07557_),
    .Y(_07732_));
 sky130_fd_sc_hd__o21ai_2 _30281_ (.A1(_07574_),
    .A2(_07732_),
    .B1(_07559_),
    .Y(_07733_));
 sky130_fd_sc_hd__a21oi_2 _30282_ (.A1(_07729_),
    .A2(_07731_),
    .B1(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__a21oi_4 _30283_ (.A1(_07700_),
    .A2(_07570_),
    .B1(_07734_),
    .Y(_07735_));
 sky130_fd_sc_hd__nand3_4 _30284_ (.A(_07733_),
    .B(_07729_),
    .C(_07731_),
    .Y(_07736_));
 sky130_fd_sc_hd__and2_1 _30285_ (.A(_07574_),
    .B(_07559_),
    .X(_07737_));
 sky130_fd_sc_hd__o2bb2ai_2 _30286_ (.A1_N(_07731_),
    .A2_N(_07729_),
    .B1(_07732_),
    .B2(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand2_2 _30287_ (.A(_07570_),
    .B(_07700_),
    .Y(_07739_));
 sky130_fd_sc_hd__a21oi_4 _30288_ (.A1(_07738_),
    .A2(_07736_),
    .B1(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__a21oi_4 _30289_ (.A1(_07735_),
    .A2(_07736_),
    .B1(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__nand2_1 _30290_ (.A(_07699_),
    .B(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__and3_1 _30291_ (.A(_07738_),
    .B(_07736_),
    .C(_07739_),
    .X(_07743_));
 sky130_fd_sc_hd__o211ai_4 _30292_ (.A1(_07740_),
    .A2(_07743_),
    .B1(_07692_),
    .C1(_07698_),
    .Y(_07744_));
 sky130_fd_sc_hd__nand3_4 _30293_ (.A(_07742_),
    .B(_07494_),
    .C(_07744_),
    .Y(_07745_));
 sky130_fd_sc_hd__o2bb2ai_2 _30294_ (.A1_N(_07692_),
    .A2_N(_07698_),
    .B1(_07740_),
    .B2(_07743_),
    .Y(_07746_));
 sky130_fd_sc_hd__nand3_2 _30295_ (.A(_07741_),
    .B(_07692_),
    .C(_07698_),
    .Y(_07747_));
 sky130_fd_sc_hd__nand3_4 _30296_ (.A(_07746_),
    .B(_07747_),
    .C(_07478_),
    .Y(_07748_));
 sky130_fd_sc_hd__nor2_1 _30297_ (.A(_07537_),
    .B(_07590_),
    .Y(_07749_));
 sky130_fd_sc_hd__o2bb2ai_2 _30298_ (.A1_N(_07745_),
    .A2_N(_07748_),
    .B1(_07540_),
    .B2(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__a21oi_2 _30299_ (.A1(_07470_),
    .A2(_07472_),
    .B1(_07468_),
    .Y(_07751_));
 sky130_fd_sc_hd__buf_6 _30300_ (.A(_05946_),
    .X(_07752_));
 sky130_fd_sc_hd__clkbuf_4 _30301_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07753_));
 sky130_fd_sc_hd__buf_6 _30302_ (.A(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__buf_2 _30303_ (.A(_19885_),
    .X(_07755_));
 sky130_fd_sc_hd__nand2_2 _30304_ (.A(_07754_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__a22o_2 _30305_ (.A1(_07446_),
    .A2(_05460_),
    .B1(_19886_),
    .B2(_05218_),
    .X(_07757_));
 sky130_fd_sc_hd__o21ai_1 _30306_ (.A1(_07752_),
    .A2(_07756_),
    .B1(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__nand2_2 _30307_ (.A(_19889_),
    .B(_05308_),
    .Y(_07759_));
 sky130_vsdinv _30308_ (.A(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__nand2_1 _30309_ (.A(_07758_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand2_1 _30310_ (.A(_07485_),
    .B(_07486_),
    .Y(_07762_));
 sky130_fd_sc_hd__a31oi_4 _30311_ (.A1(_07762_),
    .A2(_07479_),
    .A3(_20172_),
    .B1(_07487_),
    .Y(_07763_));
 sky130_fd_sc_hd__o211ai_4 _30312_ (.A1(_07752_),
    .A2(_07756_),
    .B1(_07759_),
    .C1(_07757_),
    .Y(_07764_));
 sky130_fd_sc_hd__nand3_4 _30313_ (.A(_07761_),
    .B(_07763_),
    .C(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__nand2_1 _30314_ (.A(_07758_),
    .B(_07759_),
    .Y(_07766_));
 sky130_fd_sc_hd__nor2_2 _30315_ (.A(_07752_),
    .B(_07756_),
    .Y(_07767_));
 sky130_fd_sc_hd__nand3b_2 _30316_ (.A_N(_07767_),
    .B(_07760_),
    .C(_07757_),
    .Y(_07768_));
 sky130_fd_sc_hd__o21bai_2 _30317_ (.A1(_07480_),
    .A2(_07484_),
    .B1_N(_07487_),
    .Y(_07769_));
 sky130_fd_sc_hd__nand3_4 _30318_ (.A(_07766_),
    .B(_07768_),
    .C(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__nor2_4 _30319_ (.A(_07452_),
    .B(_07448_),
    .Y(_07771_));
 sky130_fd_sc_hd__o2bb2ai_4 _30320_ (.A1_N(_07765_),
    .A2_N(_07770_),
    .B1(_07454_),
    .B2(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__nor2_4 _30321_ (.A(_07454_),
    .B(_07771_),
    .Y(_07773_));
 sky130_fd_sc_hd__nand3_4 _30322_ (.A(_07770_),
    .B(_07765_),
    .C(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__nand2_4 _30323_ (.A(_07466_),
    .B(_07456_),
    .Y(_07775_));
 sky130_fd_sc_hd__a21oi_4 _30324_ (.A1(_07772_),
    .A2(_07774_),
    .B1(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__nand2_2 _30325_ (.A(_07765_),
    .B(_07773_),
    .Y(_07777_));
 sky130_vsdinv _30326_ (.A(_07770_),
    .Y(_07778_));
 sky130_fd_sc_hd__o211a_1 _30327_ (.A1(_07777_),
    .A2(_07778_),
    .B1(_07775_),
    .C1(_07772_),
    .X(_07779_));
 sky130_fd_sc_hd__o21ai_4 _30328_ (.A1(_07419_),
    .A2(_07416_),
    .B1(_07423_),
    .Y(_07780_));
 sky130_fd_sc_hd__nand2_2 _30329_ (.A(_06543_),
    .B(_20155_),
    .Y(_07781_));
 sky130_fd_sc_hd__nand2_4 _30330_ (.A(_19895_),
    .B(_20151_),
    .Y(_07782_));
 sky130_fd_sc_hd__nor2_4 _30331_ (.A(_07781_),
    .B(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__and2_1 _30332_ (.A(_07781_),
    .B(_07782_),
    .X(_07784_));
 sky130_fd_sc_hd__buf_4 _30333_ (.A(\pcpi_mul.rs2[12] ),
    .X(_07785_));
 sky130_fd_sc_hd__nand2_2 _30334_ (.A(_07785_),
    .B(_05689_),
    .Y(_07786_));
 sky130_fd_sc_hd__o21bai_2 _30335_ (.A1(_07783_),
    .A2(_07784_),
    .B1_N(_07786_),
    .Y(_07787_));
 sky130_fd_sc_hd__or2_1 _30336_ (.A(_07781_),
    .B(_07782_),
    .X(_07788_));
 sky130_fd_sc_hd__nand2_1 _30337_ (.A(_07781_),
    .B(_07782_),
    .Y(_07789_));
 sky130_fd_sc_hd__nand3_2 _30338_ (.A(_07788_),
    .B(_07789_),
    .C(_07786_),
    .Y(_07790_));
 sky130_fd_sc_hd__nand3b_4 _30339_ (.A_N(_07780_),
    .B(_07787_),
    .C(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__o21ai_2 _30340_ (.A1(_07783_),
    .A2(_07784_),
    .B1(_07786_),
    .Y(_07792_));
 sky130_fd_sc_hd__a21oi_2 _30341_ (.A1(_07781_),
    .A2(_07782_),
    .B1(_07786_),
    .Y(_07793_));
 sky130_fd_sc_hd__nand2_1 _30342_ (.A(_07788_),
    .B(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__nand3_4 _30343_ (.A(_07792_),
    .B(_07794_),
    .C(_07780_),
    .Y(_07795_));
 sky130_fd_sc_hd__and4_2 _30344_ (.A(_06627_),
    .B(_06106_),
    .C(_06695_),
    .D(_06841_),
    .X(_07796_));
 sky130_fd_sc_hd__a22o_1 _30345_ (.A1(_06627_),
    .A2(_05826_),
    .B1(_06534_),
    .B2(_07024_),
    .X(_07797_));
 sky130_fd_sc_hd__nand2_1 _30346_ (.A(_19908_),
    .B(_07028_),
    .Y(_07798_));
 sky130_vsdinv _30347_ (.A(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__nand2_1 _30348_ (.A(_07797_),
    .B(_07799_),
    .Y(_07800_));
 sky130_fd_sc_hd__a22oi_4 _30349_ (.A1(_06344_),
    .A2(_07033_),
    .B1(_06909_),
    .B2(_05999_),
    .Y(_07801_));
 sky130_fd_sc_hd__o21ai_1 _30350_ (.A1(_07801_),
    .A2(_07796_),
    .B1(_07798_),
    .Y(_07802_));
 sky130_fd_sc_hd__o21ai_1 _30351_ (.A1(_07796_),
    .A2(_07800_),
    .B1(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__a21o_1 _30352_ (.A1(_07791_),
    .A2(_07795_),
    .B1(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__nand3_1 _30353_ (.A(_07791_),
    .B(_07795_),
    .C(_07803_),
    .Y(_07805_));
 sky130_fd_sc_hd__nand2_2 _30354_ (.A(_07804_),
    .B(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__o21ai_2 _30355_ (.A1(_07776_),
    .A2(_07779_),
    .B1(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__a21o_1 _30356_ (.A1(_07772_),
    .A2(_07774_),
    .B1(_07775_),
    .X(_07808_));
 sky130_fd_sc_hd__nand3_4 _30357_ (.A(_07772_),
    .B(_07775_),
    .C(_07774_),
    .Y(_07809_));
 sky130_fd_sc_hd__o21a_2 _30358_ (.A1(_07796_),
    .A2(_07800_),
    .B1(_07802_),
    .X(_07810_));
 sky130_fd_sc_hd__a21o_1 _30359_ (.A1(_07791_),
    .A2(_07795_),
    .B1(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__nand3_1 _30360_ (.A(_07791_),
    .B(_07810_),
    .C(_07795_),
    .Y(_07812_));
 sky130_fd_sc_hd__nand2_2 _30361_ (.A(_07811_),
    .B(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__nand3_2 _30362_ (.A(_07808_),
    .B(_07809_),
    .C(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__nand3_4 _30363_ (.A(_07751_),
    .B(_07807_),
    .C(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__o21ai_2 _30364_ (.A1(_07776_),
    .A2(_07779_),
    .B1(_07813_),
    .Y(_07816_));
 sky130_fd_sc_hd__a21o_1 _30365_ (.A1(_07428_),
    .A2(_07432_),
    .B1(_07442_),
    .X(_07817_));
 sky130_fd_sc_hd__nand2_1 _30366_ (.A(_07817_),
    .B(_07443_),
    .Y(_07818_));
 sky130_fd_sc_hd__o21ai_2 _30367_ (.A1(_07818_),
    .A2(_07465_),
    .B1(_07471_),
    .Y(_07819_));
 sky130_fd_sc_hd__nand3_2 _30368_ (.A(_07808_),
    .B(_07809_),
    .C(_07806_),
    .Y(_07820_));
 sky130_fd_sc_hd__nand3_4 _30369_ (.A(_07816_),
    .B(_07819_),
    .C(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__inv_8 _30370_ (.A(_19865_),
    .Y(_07822_));
 sky130_fd_sc_hd__nor2_8 _30371_ (.A(_07822_),
    .B(_04839_),
    .Y(_07823_));
 sky130_vsdinv _30372_ (.A(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__nand2_2 _30373_ (.A(\pcpi_mul.rs2[20] ),
    .B(\pcpi_mul.rs1[1] ),
    .Y(_07825_));
 sky130_fd_sc_hd__nand3b_4 _30374_ (.A_N(_07825_),
    .B(_19873_),
    .C(_05313_),
    .Y(_07826_));
 sky130_fd_sc_hd__buf_4 _30375_ (.A(\pcpi_mul.rs2[19] ),
    .X(_07827_));
 sky130_fd_sc_hd__nand2_1 _30376_ (.A(_07827_),
    .B(_05299_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_2 _30377_ (.A(_07825_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand2_2 _30378_ (.A(_19876_),
    .B(_05176_),
    .Y(_07830_));
 sky130_fd_sc_hd__a21o_1 _30379_ (.A1(_07826_),
    .A2(_07829_),
    .B1(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__nand3_1 _30380_ (.A(_07826_),
    .B(_07830_),
    .C(_07829_),
    .Y(_07832_));
 sky130_fd_sc_hd__nand2_2 _30381_ (.A(_07831_),
    .B(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__nor2_1 _30382_ (.A(_07824_),
    .B(_07833_),
    .Y(_07834_));
 sky130_vsdinv _30383_ (.A(_07833_),
    .Y(_07835_));
 sky130_fd_sc_hd__nor2_1 _30384_ (.A(_07823_),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__nor2_1 _30385_ (.A(_07834_),
    .B(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__a21boi_2 _30386_ (.A1(_07815_),
    .A2(_07821_),
    .B1_N(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__o211a_2 _30387_ (.A1(_07834_),
    .A2(_07836_),
    .B1(_07821_),
    .C1(_07815_),
    .X(_07839_));
 sky130_fd_sc_hd__o22ai_4 _30388_ (.A1(_07489_),
    .A2(_07603_),
    .B1(_07838_),
    .B2(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__nand3b_4 _30389_ (.A_N(_07837_),
    .B(_07815_),
    .C(_07821_),
    .Y(_07841_));
 sky130_fd_sc_hd__nor2_2 _30390_ (.A(_07489_),
    .B(_07475_),
    .Y(_07842_));
 sky130_fd_sc_hd__nor2_8 _30391_ (.A(_07824_),
    .B(_07835_),
    .Y(_07843_));
 sky130_fd_sc_hd__nor2_1 _30392_ (.A(_07823_),
    .B(_07833_),
    .Y(_07844_));
 sky130_fd_sc_hd__o2bb2ai_2 _30393_ (.A1_N(_07821_),
    .A2_N(_07815_),
    .B1(_07843_),
    .B2(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__o2111ai_4 _30394_ (.A1(_07492_),
    .A2(_07491_),
    .B1(_07841_),
    .C1(_07842_),
    .D1(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__nand2_2 _30395_ (.A(_07840_),
    .B(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand2_4 _30396_ (.A(_07597_),
    .B(_07591_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand3b_4 _30397_ (.A_N(_07848_),
    .B(_07745_),
    .C(_07748_),
    .Y(_07849_));
 sky130_fd_sc_hd__nand3_4 _30398_ (.A(_07750_),
    .B(_07847_),
    .C(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__a21o_1 _30399_ (.A1(_07750_),
    .A2(_07849_),
    .B1(_07847_),
    .X(_07851_));
 sky130_fd_sc_hd__nand3_4 _30400_ (.A(_07657_),
    .B(_07850_),
    .C(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__a21oi_4 _30401_ (.A1(_07745_),
    .A2(_07748_),
    .B1(_07848_),
    .Y(_07853_));
 sky130_fd_sc_hd__nand3_4 _30402_ (.A(_07745_),
    .B(_07748_),
    .C(_07848_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand3_4 _30403_ (.A(_07854_),
    .B(_07840_),
    .C(_07846_),
    .Y(_07855_));
 sky130_fd_sc_hd__o21ai_4 _30404_ (.A1(_07853_),
    .A2(_07855_),
    .B1(_07850_),
    .Y(_07856_));
 sky130_fd_sc_hd__nand3_4 _30405_ (.A(_07856_),
    .B(_07498_),
    .C(_07608_),
    .Y(_07857_));
 sky130_fd_sc_hd__nand2_1 _30406_ (.A(_07593_),
    .B(_07599_),
    .Y(_07858_));
 sky130_fd_sc_hd__and2_1 _30407_ (.A(_07858_),
    .B(_07598_),
    .X(_07859_));
 sky130_vsdinv _30408_ (.A(_07577_),
    .Y(_07860_));
 sky130_fd_sc_hd__nand2_4 _30409_ (.A(_07860_),
    .B(_07581_),
    .Y(_07861_));
 sky130_vsdinv _30410_ (.A(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__nand2_1 _30411_ (.A(_07859_),
    .B(_07862_),
    .Y(_07863_));
 sky130_fd_sc_hd__nand2_2 _30412_ (.A(_07858_),
    .B(_07598_),
    .Y(_07864_));
 sky130_fd_sc_hd__nand2_2 _30413_ (.A(_07864_),
    .B(_07861_),
    .Y(_07865_));
 sky130_fd_sc_hd__nand2_2 _30414_ (.A(_07863_),
    .B(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__nand3_2 _30415_ (.A(_07852_),
    .B(_07857_),
    .C(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__a21o_1 _30416_ (.A1(_07852_),
    .A2(_07857_),
    .B1(_07866_),
    .X(_07868_));
 sky130_fd_sc_hd__o2111ai_4 _30417_ (.A1(_07655_),
    .A2(_07620_),
    .B1(_07618_),
    .C1(_07867_),
    .D1(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__o21ai_2 _30418_ (.A1(_07655_),
    .A2(_07620_),
    .B1(_07618_),
    .Y(_07870_));
 sky130_vsdinv _30419_ (.A(_07865_),
    .Y(_07871_));
 sky130_vsdinv _30420_ (.A(_07863_),
    .Y(_07872_));
 sky130_fd_sc_hd__o2bb2ai_2 _30421_ (.A1_N(_07857_),
    .A2_N(_07852_),
    .B1(_07871_),
    .B2(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__xor2_4 _30422_ (.A(_07861_),
    .B(_07864_),
    .X(_07874_));
 sky130_fd_sc_hd__nand3_4 _30423_ (.A(_07874_),
    .B(_07852_),
    .C(_07857_),
    .Y(_07875_));
 sky130_fd_sc_hd__nand3_4 _30424_ (.A(_07870_),
    .B(_07873_),
    .C(_07875_),
    .Y(_07876_));
 sky130_fd_sc_hd__nand2_1 _30425_ (.A(_07869_),
    .B(_07876_),
    .Y(_07877_));
 sky130_vsdinv _30426_ (.A(_07616_),
    .Y(_07878_));
 sky130_fd_sc_hd__a22oi_4 _30427_ (.A1(_07877_),
    .A2(_07878_),
    .B1(_07630_),
    .B2(_07641_),
    .Y(_07879_));
 sky130_fd_sc_hd__nand3_4 _30428_ (.A(_07869_),
    .B(_07616_),
    .C(_07876_),
    .Y(_07880_));
 sky130_fd_sc_hd__o2bb2ai_2 _30429_ (.A1_N(_07869_),
    .A2_N(_07876_),
    .B1(_07612_),
    .B2(_07615_),
    .Y(_07881_));
 sky130_fd_sc_hd__o21ai_2 _30430_ (.A1(_07385_),
    .A2(_07635_),
    .B1(_07641_),
    .Y(_07882_));
 sky130_fd_sc_hd__a21oi_4 _30431_ (.A1(_07881_),
    .A2(_07880_),
    .B1(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__a21oi_4 _30432_ (.A1(_07879_),
    .A2(_07880_),
    .B1(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__a21oi_1 _30433_ (.A1(_07654_),
    .A2(_07643_),
    .B1(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__and3_1 _30434_ (.A(_07654_),
    .B(_07643_),
    .C(_07884_),
    .X(_07886_));
 sky130_fd_sc_hd__nor2_1 _30435_ (.A(_07885_),
    .B(_07886_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _30436_ (.A(_07852_),
    .B(_07866_),
    .Y(_07887_));
 sky130_fd_sc_hd__and2b_1 _30437_ (.A_N(_07735_),
    .B(_07736_),
    .X(_07888_));
 sky130_fd_sc_hd__a21oi_4 _30438_ (.A1(_07854_),
    .A2(_07748_),
    .B1(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__and3_2 _30439_ (.A(_07854_),
    .B(_07748_),
    .C(_07888_),
    .X(_07890_));
 sky130_fd_sc_hd__a22oi_4 _30440_ (.A1(_07446_),
    .A2(_05218_),
    .B1(_06637_),
    .B2(_05389_),
    .Y(_07891_));
 sky130_fd_sc_hd__and4_4 _30441_ (.A(_07754_),
    .B(_07755_),
    .C(_20158_),
    .D(_05289_),
    .X(_07892_));
 sky130_fd_sc_hd__buf_4 _30442_ (.A(\pcpi_mul.rs2[15] ),
    .X(_07893_));
 sky130_fd_sc_hd__nand2_2 _30443_ (.A(_07893_),
    .B(_20155_),
    .Y(_07894_));
 sky130_fd_sc_hd__o21ai_2 _30444_ (.A1(_07891_),
    .A2(_07892_),
    .B1(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_1 _30445_ (.A(_06927_),
    .B(_05480_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand3b_4 _30446_ (.A_N(_07896_),
    .B(_07449_),
    .C(_05684_),
    .Y(_07897_));
 sky130_vsdinv _30447_ (.A(_07894_),
    .Y(_07898_));
 sky130_fd_sc_hd__a22o_4 _30448_ (.A1(_07446_),
    .A2(_05392_),
    .B1(_19886_),
    .B2(_07417_),
    .X(_07899_));
 sky130_fd_sc_hd__nand3_4 _30449_ (.A(_07897_),
    .B(_07898_),
    .C(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__buf_6 _30450_ (.A(_20173_),
    .X(_07901_));
 sky130_fd_sc_hd__buf_6 _30451_ (.A(_07827_),
    .X(_07902_));
 sky130_fd_sc_hd__a22oi_4 _30452_ (.A1(_19870_),
    .A2(_07901_),
    .B1(_07902_),
    .B2(_05179_),
    .Y(_07903_));
 sky130_fd_sc_hd__o21ai_4 _30453_ (.A1(_07830_),
    .A2(_07903_),
    .B1(_07826_),
    .Y(_07904_));
 sky130_fd_sc_hd__nand3_4 _30454_ (.A(_07895_),
    .B(_07900_),
    .C(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__o21ai_2 _30455_ (.A1(_07891_),
    .A2(_07892_),
    .B1(_07898_),
    .Y(_07906_));
 sky130_fd_sc_hd__nand3_4 _30456_ (.A(_07897_),
    .B(_07894_),
    .C(_07899_),
    .Y(_07907_));
 sky130_fd_sc_hd__o21ai_2 _30457_ (.A1(_07825_),
    .A2(_07828_),
    .B1(_07830_),
    .Y(_07908_));
 sky130_fd_sc_hd__nand2_4 _30458_ (.A(_07908_),
    .B(_07829_),
    .Y(_07909_));
 sky130_fd_sc_hd__nand3_2 _30459_ (.A(_07906_),
    .B(_07907_),
    .C(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__a21oi_4 _30460_ (.A1(_07757_),
    .A2(_07760_),
    .B1(_07767_),
    .Y(_07911_));
 sky130_vsdinv _30461_ (.A(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__a21o_2 _30462_ (.A1(_07905_),
    .A2(_07910_),
    .B1(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__a31oi_4 _30463_ (.A1(_07906_),
    .A2(_07907_),
    .A3(_07909_),
    .B1(_07911_),
    .Y(_07914_));
 sky130_fd_sc_hd__nand2_4 _30464_ (.A(_07914_),
    .B(_07905_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_4 _30465_ (.A(_07777_),
    .B(_07770_),
    .Y(_07916_));
 sky130_fd_sc_hd__a21oi_4 _30466_ (.A1(_07913_),
    .A2(_07915_),
    .B1(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__and3_1 _30467_ (.A(_07895_),
    .B(_07900_),
    .C(_07904_),
    .X(_07918_));
 sky130_fd_sc_hd__nand2_1 _30468_ (.A(_07910_),
    .B(_07912_),
    .Y(_07919_));
 sky130_fd_sc_hd__o211a_1 _30469_ (.A1(_07918_),
    .A2(_07919_),
    .B1(_07913_),
    .C1(_07916_),
    .X(_07920_));
 sky130_fd_sc_hd__nor2_2 _30470_ (.A(_07783_),
    .B(_07793_),
    .Y(_07921_));
 sky130_fd_sc_hd__buf_6 _30471_ (.A(_06356_),
    .X(_07922_));
 sky130_fd_sc_hd__a22oi_4 _30472_ (.A1(_07922_),
    .A2(_05571_),
    .B1(_06207_),
    .B2(_05827_),
    .Y(_07923_));
 sky130_fd_sc_hd__nand2_2 _30473_ (.A(_06356_),
    .B(_05453_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_2 _30474_ (.A(_19895_),
    .B(_20148_),
    .Y(_07925_));
 sky130_fd_sc_hd__nor2_4 _30475_ (.A(_07924_),
    .B(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nand2_2 _30476_ (.A(_07785_),
    .B(_05670_),
    .Y(_07927_));
 sky130_vsdinv _30477_ (.A(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__o21ai_2 _30478_ (.A1(_07923_),
    .A2(_07926_),
    .B1(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand3b_2 _30479_ (.A_N(_07924_),
    .B(_19896_),
    .C(_06289_),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_2 _30480_ (.A(_07924_),
    .B(_07925_),
    .Y(_07931_));
 sky130_fd_sc_hd__nand3_4 _30481_ (.A(_07930_),
    .B(_07927_),
    .C(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__nand3_4 _30482_ (.A(_07921_),
    .B(_07929_),
    .C(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__a22oi_4 _30483_ (.A1(_06630_),
    .A2(_20142_),
    .B1(_06631_),
    .B2(_20138_),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_1 _30484_ (.A(_06622_),
    .B(_20141_),
    .Y(_07935_));
 sky130_fd_sc_hd__nand2_1 _30485_ (.A(_06044_),
    .B(_07028_),
    .Y(_07936_));
 sky130_fd_sc_hd__nor2_1 _30486_ (.A(_07935_),
    .B(_07936_),
    .Y(_07937_));
 sky130_fd_sc_hd__nand2_2 _30487_ (.A(_06051_),
    .B(_07661_),
    .Y(_07938_));
 sky130_fd_sc_hd__o21bai_1 _30488_ (.A1(_07934_),
    .A2(_07937_),
    .B1_N(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand3b_2 _30489_ (.A_N(_07935_),
    .B(_05657_),
    .C(_07185_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand2_1 _30490_ (.A(_07935_),
    .B(_07936_),
    .Y(_07941_));
 sky130_fd_sc_hd__nand3_1 _30491_ (.A(_07940_),
    .B(_07941_),
    .C(_07938_),
    .Y(_07942_));
 sky130_fd_sc_hd__nand2_2 _30492_ (.A(_07939_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_2 _30493_ (.A(_07933_),
    .B(_07943_),
    .Y(_07944_));
 sky130_fd_sc_hd__a21o_1 _30494_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_07921_),
    .X(_07945_));
 sky130_vsdinv _30495_ (.A(_07945_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand2_1 _30496_ (.A(_07945_),
    .B(_07933_),
    .Y(_07947_));
 sky130_vsdinv _30497_ (.A(_07943_),
    .Y(_07948_));
 sky130_fd_sc_hd__nand2_1 _30498_ (.A(_07947_),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__o21ai_4 _30499_ (.A1(_07944_),
    .A2(_07946_),
    .B1(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__o21ai_2 _30500_ (.A1(_07917_),
    .A2(_07920_),
    .B1(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__o21ai_2 _30501_ (.A1(_07813_),
    .A2(_07776_),
    .B1(_07809_),
    .Y(_07952_));
 sky130_fd_sc_hd__a21o_1 _30502_ (.A1(_07913_),
    .A2(_07915_),
    .B1(_07916_),
    .X(_07953_));
 sky130_fd_sc_hd__nand3_4 _30503_ (.A(_07916_),
    .B(_07913_),
    .C(_07915_),
    .Y(_07954_));
 sky130_fd_sc_hd__nand2_1 _30504_ (.A(_07947_),
    .B(_07943_),
    .Y(_07955_));
 sky130_fd_sc_hd__nand3_1 _30505_ (.A(_07948_),
    .B(_07945_),
    .C(_07933_),
    .Y(_07956_));
 sky130_fd_sc_hd__nand2_1 _30506_ (.A(_07955_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__nand3_2 _30507_ (.A(_07953_),
    .B(_07954_),
    .C(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__nand3_4 _30508_ (.A(_07951_),
    .B(_07952_),
    .C(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__o21ai_2 _30509_ (.A1(_07917_),
    .A2(_07920_),
    .B1(_07957_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand2_1 _30510_ (.A(_07813_),
    .B(_07809_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2_1 _30511_ (.A(_07961_),
    .B(_07808_),
    .Y(_07962_));
 sky130_fd_sc_hd__nand3_2 _30512_ (.A(_07953_),
    .B(_07954_),
    .C(_07950_),
    .Y(_07963_));
 sky130_fd_sc_hd__nand3_4 _30513_ (.A(_07960_),
    .B(_07962_),
    .C(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__clkbuf_8 _30514_ (.A(_19862_),
    .X(_07965_));
 sky130_fd_sc_hd__nand2_2 _30515_ (.A(_07965_),
    .B(_05214_),
    .Y(_07966_));
 sky130_fd_sc_hd__buf_8 _30516_ (.A(_19865_),
    .X(_07967_));
 sky130_fd_sc_hd__nand2_2 _30517_ (.A(_07967_),
    .B(_05146_),
    .Y(_07968_));
 sky130_fd_sc_hd__nand2_1 _30518_ (.A(_07966_),
    .B(_07968_),
    .Y(_07969_));
 sky130_fd_sc_hd__nor2_4 _30519_ (.A(_07966_),
    .B(_07968_),
    .Y(_07970_));
 sky130_vsdinv _30520_ (.A(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__nand2_2 _30521_ (.A(_19869_),
    .B(_05299_),
    .Y(_07972_));
 sky130_fd_sc_hd__buf_8 _30522_ (.A(_19872_),
    .X(_07973_));
 sky130_fd_sc_hd__nand3b_4 _30523_ (.A_N(_07972_),
    .B(_07973_),
    .C(_05245_),
    .Y(_07974_));
 sky130_fd_sc_hd__nand2_2 _30524_ (.A(_07827_),
    .B(_05602_),
    .Y(_07975_));
 sky130_fd_sc_hd__nand2_4 _30525_ (.A(_07972_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__a22o_1 _30526_ (.A1(_19878_),
    .A2(_20166_),
    .B1(_07974_),
    .B2(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__nand2_2 _30527_ (.A(_19876_),
    .B(_05549_),
    .Y(_07978_));
 sky130_fd_sc_hd__nand3b_4 _30528_ (.A_N(_07978_),
    .B(_07974_),
    .C(_07976_),
    .Y(_07979_));
 sky130_fd_sc_hd__a22o_4 _30529_ (.A1(_07969_),
    .A2(_07971_),
    .B1(_07977_),
    .B2(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__nand2_1 _30530_ (.A(_07971_),
    .B(_07969_),
    .Y(_07981_));
 sky130_fd_sc_hd__nand3b_4 _30531_ (.A_N(_07981_),
    .B(_07977_),
    .C(_07979_),
    .Y(_07982_));
 sky130_fd_sc_hd__a21oi_4 _30532_ (.A1(_07980_),
    .A2(_07982_),
    .B1(_07843_),
    .Y(_07983_));
 sky130_fd_sc_hd__nand3_4 _30533_ (.A(_07843_),
    .B(_07980_),
    .C(_07982_),
    .Y(_07984_));
 sky130_vsdinv _30534_ (.A(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__o2bb2ai_2 _30535_ (.A1_N(_07959_),
    .A2_N(_07964_),
    .B1(_07983_),
    .B2(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__nor2_2 _30536_ (.A(_07983_),
    .B(_07985_),
    .Y(_07987_));
 sky130_fd_sc_hd__nand3_4 _30537_ (.A(_07959_),
    .B(_07964_),
    .C(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__a21oi_4 _30538_ (.A1(_07986_),
    .A2(_07988_),
    .B1(_07839_),
    .Y(_07989_));
 sky130_fd_sc_hd__nand2_2 _30539_ (.A(_07986_),
    .B(_07988_),
    .Y(_07990_));
 sky130_fd_sc_hd__nor2_4 _30540_ (.A(_07841_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__nand2_1 _30541_ (.A(_07791_),
    .B(_07810_),
    .Y(_07992_));
 sky130_fd_sc_hd__nand2_1 _30542_ (.A(_07992_),
    .B(_07795_),
    .Y(_07993_));
 sky130_fd_sc_hd__a22oi_4 _30543_ (.A1(_07660_),
    .A2(_06715_),
    .B1(_05413_),
    .B2(_06813_),
    .Y(_07994_));
 sky130_fd_sc_hd__clkinv_8 _30544_ (.A(net473),
    .Y(_07995_));
 sky130_fd_sc_hd__nand3_4 _30545_ (.A(_06659_),
    .B(_05724_),
    .C(_06294_),
    .Y(_07996_));
 sky130_fd_sc_hd__nor2_4 _30546_ (.A(_07995_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__nand2_2 _30547_ (.A(_05601_),
    .B(_06701_),
    .Y(_07998_));
 sky130_vsdinv _30548_ (.A(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__o21ai_2 _30549_ (.A1(_07994_),
    .A2(_07997_),
    .B1(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21oi_2 _30550_ (.A1(_07797_),
    .A2(_07799_),
    .B1(_07796_),
    .Y(_08001_));
 sky130_fd_sc_hd__buf_6 _30551_ (.A(_20128_),
    .X(_08002_));
 sky130_fd_sc_hd__a22o_2 _30552_ (.A1(_06478_),
    .A2(_06437_),
    .B1(_06097_),
    .B2(_08002_),
    .X(_08003_));
 sky130_fd_sc_hd__o211ai_2 _30553_ (.A1(_07995_),
    .A2(_07996_),
    .B1(_07998_),
    .C1(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__nand3_4 _30554_ (.A(_08000_),
    .B(_08001_),
    .C(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__o21ai_2 _30555_ (.A1(_07994_),
    .A2(_07997_),
    .B1(_07998_),
    .Y(_08006_));
 sky130_fd_sc_hd__nand2_1 _30556_ (.A(_19901_),
    .B(_05822_),
    .Y(_08007_));
 sky130_fd_sc_hd__buf_6 _30557_ (.A(_06153_),
    .X(_08008_));
 sky130_fd_sc_hd__nand3b_2 _30558_ (.A_N(_08007_),
    .B(_07333_),
    .C(_08008_),
    .Y(_08009_));
 sky130_fd_sc_hd__o21ai_2 _30559_ (.A1(_07798_),
    .A2(_07801_),
    .B1(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__o211ai_2 _30560_ (.A1(_07995_),
    .A2(_07996_),
    .B1(_07999_),
    .C1(_08003_),
    .Y(_08011_));
 sky130_fd_sc_hd__nand3_4 _30561_ (.A(_08006_),
    .B(_08010_),
    .C(_08011_),
    .Y(_08012_));
 sky130_fd_sc_hd__a21o_2 _30562_ (.A1(_07668_),
    .A2(_07667_),
    .B1(_07663_),
    .X(_08013_));
 sky130_fd_sc_hd__nand3_4 _30563_ (.A(_08005_),
    .B(_08012_),
    .C(_08013_),
    .Y(_08014_));
 sky130_fd_sc_hd__a21o_1 _30564_ (.A1(_08005_),
    .A2(_08012_),
    .B1(_08013_),
    .X(_08015_));
 sky130_fd_sc_hd__nand3_4 _30565_ (.A(_07993_),
    .B(_08014_),
    .C(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__a21oi_2 _30566_ (.A1(_08005_),
    .A2(_08012_),
    .B1(_08013_),
    .Y(_08017_));
 sky130_fd_sc_hd__and3_1 _30567_ (.A(_08005_),
    .B(_08012_),
    .C(_08013_),
    .X(_08018_));
 sky130_fd_sc_hd__a21boi_4 _30568_ (.A1(_07791_),
    .A2(_07810_),
    .B1_N(_07795_),
    .Y(_08019_));
 sky130_fd_sc_hd__o21ai_4 _30569_ (.A1(_08017_),
    .A2(_08018_),
    .B1(_08019_),
    .Y(_08020_));
 sky130_vsdinv _30570_ (.A(_07674_),
    .Y(_08021_));
 sky130_fd_sc_hd__nor2_1 _30571_ (.A(_07677_),
    .B(_07682_),
    .Y(_08022_));
 sky130_fd_sc_hd__o2bb2ai_2 _30572_ (.A1_N(_08016_),
    .A2_N(_08020_),
    .B1(_08021_),
    .B2(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_1 _30573_ (.A(_07683_),
    .B(_07670_),
    .Y(_08024_));
 sky130_fd_sc_hd__nand3_2 _30574_ (.A(_08020_),
    .B(_08016_),
    .C(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__o21ai_2 _30575_ (.A1(_07690_),
    .A2(_07681_),
    .B1(_07689_),
    .Y(_08026_));
 sky130_fd_sc_hd__nand3_4 _30576_ (.A(_08023_),
    .B(_08025_),
    .C(_08026_),
    .Y(_08027_));
 sky130_vsdinv _30577_ (.A(_07678_),
    .Y(_08028_));
 sky130_fd_sc_hd__o2bb2ai_1 _30578_ (.A1_N(_08016_),
    .A2_N(_08020_),
    .B1(_07682_),
    .B2(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_1 _30579_ (.A(_07689_),
    .B(_07690_),
    .Y(_08030_));
 sky130_fd_sc_hd__nand2_1 _30580_ (.A(_08030_),
    .B(_07688_),
    .Y(_08031_));
 sky130_vsdinv _30581_ (.A(_08024_),
    .Y(_08032_));
 sky130_fd_sc_hd__nand3_2 _30582_ (.A(_08020_),
    .B(_08016_),
    .C(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__nand3_4 _30583_ (.A(_08029_),
    .B(_08031_),
    .C(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand2_1 _30584_ (.A(_08027_),
    .B(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__buf_4 _30585_ (.A(\pcpi_mul.rs1[22] ),
    .X(_08036_));
 sky130_fd_sc_hd__inv_8 _30586_ (.A(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__buf_6 _30587_ (.A(_08037_),
    .X(_08038_));
 sky130_vsdinv _30588_ (.A(\pcpi_mul.rs1[17] ),
    .Y(_08039_));
 sky130_fd_sc_hd__buf_8 _30589_ (.A(_08039_),
    .X(_08040_));
 sky130_fd_sc_hd__nand3_4 _30590_ (.A(_05376_),
    .B(_05211_),
    .C(_06993_),
    .Y(_08041_));
 sky130_fd_sc_hd__buf_4 _30591_ (.A(_20117_),
    .X(_08042_));
 sky130_fd_sc_hd__a22o_2 _30592_ (.A1(_06986_),
    .A2(_07702_),
    .B1(_06988_),
    .B2(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__o21ai_2 _30593_ (.A1(_08040_),
    .A2(_08041_),
    .B1(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__o21ai_4 _30594_ (.A1(net470),
    .A2(_08038_),
    .B1(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__nor2_4 _30595_ (.A(_08040_),
    .B(_08041_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_8 _30596_ (.A(_04836_),
    .B(_08037_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand3b_4 _30597_ (.A_N(_08046_),
    .B(_08043_),
    .C(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__o21ai_4 _30598_ (.A1(_07710_),
    .A2(_07706_),
    .B1(_07704_),
    .Y(_08049_));
 sky130_fd_sc_hd__a21oi_4 _30599_ (.A1(_08045_),
    .A2(_08048_),
    .B1(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__o211a_1 _30600_ (.A1(_07711_),
    .A2(_07714_),
    .B1(_08048_),
    .C1(_08045_),
    .X(_08051_));
 sky130_fd_sc_hd__buf_6 _30601_ (.A(\pcpi_mul.rs1[21] ),
    .X(_08052_));
 sky130_fd_sc_hd__buf_4 _30602_ (.A(\pcpi_mul.rs1[20] ),
    .X(_08053_));
 sky130_fd_sc_hd__nand2_1 _30603_ (.A(_05282_),
    .B(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__a21o_1 _30604_ (.A1(_05821_),
    .A2(_08052_),
    .B1(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__buf_4 _30605_ (.A(\pcpi_mul.rs1[20] ),
    .X(_08056_));
 sky130_fd_sc_hd__buf_4 _30606_ (.A(\pcpi_mul.rs1[21] ),
    .X(_08057_));
 sky130_fd_sc_hd__nand2_1 _30607_ (.A(_05477_),
    .B(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__a21o_1 _30608_ (.A1(_06314_),
    .A2(_08056_),
    .B1(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__buf_6 _30609_ (.A(_07233_),
    .X(_08060_));
 sky130_fd_sc_hd__nand2_2 _30610_ (.A(_05830_),
    .B(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__a21o_2 _30611_ (.A1(_08055_),
    .A2(_08059_),
    .B1(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__nand3_4 _30612_ (.A(_08055_),
    .B(_08059_),
    .C(_08061_),
    .Y(_08063_));
 sky130_fd_sc_hd__nand2_4 _30613_ (.A(_08062_),
    .B(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__o21ai_2 _30614_ (.A1(_08050_),
    .A2(_08051_),
    .B1(_08064_),
    .Y(_08065_));
 sky130_fd_sc_hd__and2_1 _30615_ (.A(_08062_),
    .B(_08063_),
    .X(_08066_));
 sky130_fd_sc_hd__a21o_1 _30616_ (.A1(_08045_),
    .A2(_08048_),
    .B1(_08049_),
    .X(_08067_));
 sky130_fd_sc_hd__nand3_4 _30617_ (.A(_08045_),
    .B(_08049_),
    .C(_08048_),
    .Y(_08068_));
 sky130_fd_sc_hd__nand3_2 _30618_ (.A(_08066_),
    .B(_08067_),
    .C(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__nand2_1 _30619_ (.A(_07713_),
    .B(_07730_),
    .Y(_08070_));
 sky130_fd_sc_hd__nand2_1 _30620_ (.A(_08070_),
    .B(_07717_),
    .Y(_08071_));
 sky130_fd_sc_hd__nand3_4 _30621_ (.A(_08065_),
    .B(_08069_),
    .C(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__and2_2 _30622_ (.A(_08070_),
    .B(_07717_),
    .X(_08073_));
 sky130_fd_sc_hd__o21ai_4 _30623_ (.A1(_08050_),
    .A2(_08051_),
    .B1(_08066_),
    .Y(_08074_));
 sky130_fd_sc_hd__nand3_4 _30624_ (.A(_08067_),
    .B(_08064_),
    .C(_08068_),
    .Y(_08075_));
 sky130_fd_sc_hd__o21ba_4 _30625_ (.A1(_07721_),
    .A2(_07719_),
    .B1_N(_07728_),
    .X(_08076_));
 sky130_fd_sc_hd__a31oi_4 _30626_ (.A1(_08073_),
    .A2(_08074_),
    .A3(_08075_),
    .B1(_08076_),
    .Y(_08077_));
 sky130_fd_sc_hd__nand3_4 _30627_ (.A(_08073_),
    .B(_08074_),
    .C(_08075_),
    .Y(_08078_));
 sky130_fd_sc_hd__a21boi_4 _30628_ (.A1(_08078_),
    .A2(_08072_),
    .B1_N(_08076_),
    .Y(_08079_));
 sky130_fd_sc_hd__a21oi_4 _30629_ (.A1(_08072_),
    .A2(_08077_),
    .B1(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__nand2_1 _30630_ (.A(_08035_),
    .B(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__nand2_1 _30631_ (.A(_08078_),
    .B(_08072_),
    .Y(_08082_));
 sky130_fd_sc_hd__nor2_4 _30632_ (.A(_08076_),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__o211ai_4 _30633_ (.A1(_08079_),
    .A2(_08083_),
    .B1(_08027_),
    .C1(_08034_),
    .Y(_08084_));
 sky130_fd_sc_hd__nand3_4 _30634_ (.A(_08081_),
    .B(_07821_),
    .C(_08084_),
    .Y(_08085_));
 sky130_fd_sc_hd__o2bb2ai_2 _30635_ (.A1_N(_08027_),
    .A2_N(_08034_),
    .B1(_08083_),
    .B2(_08079_),
    .Y(_08086_));
 sky130_fd_sc_hd__nand3_2 _30636_ (.A(_08080_),
    .B(_08027_),
    .C(_08034_),
    .Y(_08087_));
 sky130_vsdinv _30637_ (.A(_07821_),
    .Y(_08088_));
 sky130_fd_sc_hd__nand3_4 _30638_ (.A(_08086_),
    .B(_08087_),
    .C(_08088_),
    .Y(_08089_));
 sky130_vsdinv _30639_ (.A(_07698_),
    .Y(_08090_));
 sky130_fd_sc_hd__a21o_2 _30640_ (.A1(_07741_),
    .A2(_07692_),
    .B1(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__a21oi_4 _30641_ (.A1(_08085_),
    .A2(_08089_),
    .B1(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__and2_1 _30642_ (.A(_07741_),
    .B(_07692_),
    .X(_08093_));
 sky130_fd_sc_hd__o211a_1 _30643_ (.A1(_08090_),
    .A2(_08093_),
    .B1(_08089_),
    .C1(_08085_),
    .X(_08094_));
 sky130_fd_sc_hd__o22ai_4 _30644_ (.A1(_07989_),
    .A2(_07991_),
    .B1(_08092_),
    .B2(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__a21o_1 _30645_ (.A1(_08085_),
    .A2(_08089_),
    .B1(_08091_),
    .X(_08096_));
 sky130_fd_sc_hd__nand2_2 _30646_ (.A(_07964_),
    .B(_07959_),
    .Y(_08097_));
 sky130_vsdinv _30647_ (.A(_07987_),
    .Y(_08098_));
 sky130_fd_sc_hd__a21oi_2 _30648_ (.A1(_08097_),
    .A2(_08098_),
    .B1(_07841_),
    .Y(_08099_));
 sky130_fd_sc_hd__a21oi_2 _30649_ (.A1(_08099_),
    .A2(_07988_),
    .B1(_07989_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand3_4 _30650_ (.A(_08085_),
    .B(_08089_),
    .C(_08091_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand3_4 _30651_ (.A(_08096_),
    .B(_08100_),
    .C(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__nand2_1 _30652_ (.A(_07845_),
    .B(_07841_),
    .Y(_08103_));
 sky130_fd_sc_hd__o22ai_4 _30653_ (.A1(_07495_),
    .A2(_08103_),
    .B1(_07853_),
    .B2(_07855_),
    .Y(_08104_));
 sky130_fd_sc_hd__a21oi_4 _30654_ (.A1(_08095_),
    .A2(_08102_),
    .B1(_08104_),
    .Y(_08105_));
 sky130_fd_sc_hd__nand2_2 _30655_ (.A(_07990_),
    .B(_07841_),
    .Y(_08106_));
 sky130_fd_sc_hd__nand2_1 _30656_ (.A(_08099_),
    .B(_07988_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand3_2 _30657_ (.A(_08101_),
    .B(_08106_),
    .C(_08107_),
    .Y(_08108_));
 sky130_fd_sc_hd__o211a_2 _30658_ (.A1(_08092_),
    .A2(_08108_),
    .B1(_08095_),
    .C1(_08104_),
    .X(_08109_));
 sky130_fd_sc_hd__o22ai_4 _30659_ (.A1(_07889_),
    .A2(_07890_),
    .B1(_08105_),
    .B2(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__a21o_1 _30660_ (.A1(_08095_),
    .A2(_08102_),
    .B1(_08104_),
    .X(_08111_));
 sky130_fd_sc_hd__nand3_4 _30661_ (.A(_08104_),
    .B(_08095_),
    .C(_08102_),
    .Y(_08112_));
 sky130_fd_sc_hd__nor2_8 _30662_ (.A(_07889_),
    .B(_07890_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand3_4 _30663_ (.A(_08111_),
    .B(_08112_),
    .C(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__a22oi_4 _30664_ (.A1(_07857_),
    .A2(_07887_),
    .B1(_08110_),
    .B2(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__o21a_1 _30665_ (.A1(_07600_),
    .A2(_07622_),
    .B1(_07498_),
    .X(_08116_));
 sky130_fd_sc_hd__nor2_1 _30666_ (.A(_07856_),
    .B(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__a21oi_1 _30667_ (.A1(_08116_),
    .A2(_07856_),
    .B1(_07866_),
    .Y(_08118_));
 sky130_fd_sc_hd__o211a_1 _30668_ (.A1(_08117_),
    .A2(_08118_),
    .B1(_08114_),
    .C1(_08110_),
    .X(_08119_));
 sky130_fd_sc_hd__o21ai_1 _30669_ (.A1(_08115_),
    .A2(_08119_),
    .B1(_07871_),
    .Y(_08120_));
 sky130_fd_sc_hd__a21boi_4 _30670_ (.A1(_07869_),
    .A2(_07616_),
    .B1_N(_07876_),
    .Y(_08121_));
 sky130_fd_sc_hd__nand2_1 _30671_ (.A(_07874_),
    .B(_07857_),
    .Y(_08122_));
 sky130_fd_sc_hd__nand2_2 _30672_ (.A(_08122_),
    .B(_07852_),
    .Y(_08123_));
 sky130_fd_sc_hd__a21o_2 _30673_ (.A1(_08110_),
    .A2(_08114_),
    .B1(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__nand3_4 _30674_ (.A(_08123_),
    .B(_08110_),
    .C(_08114_),
    .Y(_08125_));
 sky130_fd_sc_hd__nand3_2 _30675_ (.A(_08124_),
    .B(_07865_),
    .C(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__nand3_2 _30676_ (.A(_08120_),
    .B(_08121_),
    .C(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__o22ai_4 _30677_ (.A1(_07862_),
    .A2(_07859_),
    .B1(_08115_),
    .B2(_08119_),
    .Y(_08128_));
 sky130_fd_sc_hd__a21oi_1 _30678_ (.A1(_07873_),
    .A2(_07875_),
    .B1(_07870_),
    .Y(_08129_));
 sky130_fd_sc_hd__o21ai_2 _30679_ (.A1(_07878_),
    .A2(_08129_),
    .B1(_07876_),
    .Y(_08130_));
 sky130_fd_sc_hd__nand3_4 _30680_ (.A(_08124_),
    .B(_07871_),
    .C(_08125_),
    .Y(_08131_));
 sky130_fd_sc_hd__nand3_4 _30681_ (.A(_08128_),
    .B(_08130_),
    .C(_08131_),
    .Y(_08132_));
 sky130_fd_sc_hd__nand2_1 _30682_ (.A(_08127_),
    .B(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__nand2_2 _30683_ (.A(_07649_),
    .B(_07651_),
    .Y(_08134_));
 sky130_fd_sc_hd__nand3_2 _30684_ (.A(_07881_),
    .B(_07882_),
    .C(_07880_),
    .Y(_08135_));
 sky130_fd_sc_hd__a21oi_4 _30685_ (.A1(_07653_),
    .A2(_08135_),
    .B1(_07883_),
    .Y(_08136_));
 sky130_fd_sc_hd__a31oi_4 _30686_ (.A1(_08134_),
    .A2(_07644_),
    .A3(_07884_),
    .B1(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__xor2_2 _30687_ (.A(_08133_),
    .B(_08137_),
    .X(_02641_));
 sky130_fd_sc_hd__a31o_1 _30688_ (.A1(_08121_),
    .A2(_08126_),
    .A3(_08120_),
    .B1(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__nand2_2 _30689_ (.A(_08016_),
    .B(_08032_),
    .Y(_08139_));
 sky130_vsdinv _30690_ (.A(_08005_),
    .Y(_08140_));
 sky130_fd_sc_hd__and2b_1 _30691_ (.A_N(_08013_),
    .B(_08012_),
    .X(_08141_));
 sky130_fd_sc_hd__buf_4 _30692_ (.A(\pcpi_mul.rs1[16] ),
    .X(_08142_));
 sky130_fd_sc_hd__a22oi_4 _30693_ (.A1(_06095_),
    .A2(_08002_),
    .B1(_06097_),
    .B2(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand2_8 _30694_ (.A(_06701_),
    .B(_20129_),
    .Y(_08144_));
 sky130_fd_sc_hd__nor2_4 _30695_ (.A(_05860_),
    .B(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__nand2_2 _30696_ (.A(_19917_),
    .B(_07702_),
    .Y(_08146_));
 sky130_fd_sc_hd__o21ai_2 _30697_ (.A1(_08143_),
    .A2(_08145_),
    .B1(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__o21ai_2 _30698_ (.A1(_07938_),
    .A2(_07934_),
    .B1(_07940_),
    .Y(_08148_));
 sky130_fd_sc_hd__nand3_4 _30699_ (.A(_05722_),
    .B(_19914_),
    .C(_20125_),
    .Y(_08149_));
 sky130_vsdinv _30700_ (.A(_08146_),
    .Y(_08150_));
 sky130_fd_sc_hd__buf_6 _30701_ (.A(_06713_),
    .X(_08151_));
 sky130_fd_sc_hd__a22o_2 _30702_ (.A1(_06483_),
    .A2(_08151_),
    .B1(_06657_),
    .B2(_08142_),
    .X(_08152_));
 sky130_fd_sc_hd__o211ai_4 _30703_ (.A1(_07995_),
    .A2(_08149_),
    .B1(_08150_),
    .C1(_08152_),
    .Y(_08153_));
 sky130_fd_sc_hd__nand3_4 _30704_ (.A(_08147_),
    .B(_08148_),
    .C(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__o21ai_2 _30705_ (.A1(_08143_),
    .A2(_08145_),
    .B1(_08150_),
    .Y(_08155_));
 sky130_fd_sc_hd__o21ai_1 _30706_ (.A1(_07935_),
    .A2(_07936_),
    .B1(_07938_),
    .Y(_08156_));
 sky130_fd_sc_hd__nand2_1 _30707_ (.A(_08156_),
    .B(_07941_),
    .Y(_08157_));
 sky130_fd_sc_hd__o211ai_4 _30708_ (.A1(_05861_),
    .A2(_08144_),
    .B1(_08146_),
    .C1(_08152_),
    .Y(_08158_));
 sky130_fd_sc_hd__nand3_4 _30709_ (.A(_08155_),
    .B(_08157_),
    .C(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__nor2_4 _30710_ (.A(_07999_),
    .B(_07997_),
    .Y(_08160_));
 sky130_fd_sc_hd__o2bb2ai_4 _30711_ (.A1_N(_08154_),
    .A2_N(_08159_),
    .B1(_07994_),
    .B2(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__nor2_2 _30712_ (.A(_07994_),
    .B(_08160_),
    .Y(_08162_));
 sky130_fd_sc_hd__nand3_4 _30713_ (.A(_08154_),
    .B(_08159_),
    .C(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__nand2_4 _30714_ (.A(_07944_),
    .B(_07945_),
    .Y(_08164_));
 sky130_fd_sc_hd__a21oi_4 _30715_ (.A1(_08161_),
    .A2(_08163_),
    .B1(_08164_),
    .Y(_08165_));
 sky130_vsdinv _30716_ (.A(_08154_),
    .Y(_08166_));
 sky130_fd_sc_hd__nand2_1 _30717_ (.A(_08159_),
    .B(_08162_),
    .Y(_08167_));
 sky130_fd_sc_hd__o211a_1 _30718_ (.A1(_08166_),
    .A2(_08167_),
    .B1(_08161_),
    .C1(_08164_),
    .X(_08168_));
 sky130_fd_sc_hd__o22ai_4 _30719_ (.A1(_08140_),
    .A2(_08141_),
    .B1(_08165_),
    .B2(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_1 _30720_ (.A(_08005_),
    .B(_08013_),
    .Y(_08170_));
 sky130_fd_sc_hd__and2_1 _30721_ (.A(_08170_),
    .B(_08012_),
    .X(_08171_));
 sky130_fd_sc_hd__a21o_1 _30722_ (.A1(_08161_),
    .A2(_08163_),
    .B1(_08164_),
    .X(_08172_));
 sky130_fd_sc_hd__nand3_4 _30723_ (.A(_08164_),
    .B(_08161_),
    .C(_08163_),
    .Y(_08173_));
 sky130_fd_sc_hd__nand3b_4 _30724_ (.A_N(_08171_),
    .B(_08172_),
    .C(_08173_),
    .Y(_08174_));
 sky130_fd_sc_hd__a22oi_4 _30725_ (.A1(_08020_),
    .A2(_08139_),
    .B1(_08169_),
    .B2(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__nand2_2 _30726_ (.A(_08015_),
    .B(_08014_),
    .Y(_08176_));
 sky130_fd_sc_hd__nor2_2 _30727_ (.A(_08019_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__a21oi_4 _30728_ (.A1(_08176_),
    .A2(_08019_),
    .B1(_08032_),
    .Y(_08178_));
 sky130_fd_sc_hd__o211a_2 _30729_ (.A1(_08177_),
    .A2(_08178_),
    .B1(_08174_),
    .C1(_08169_),
    .X(_08179_));
 sky130_fd_sc_hd__a21o_1 _30730_ (.A1(_08047_),
    .A2(_08043_),
    .B1(_08046_),
    .X(_08180_));
 sky130_fd_sc_hd__nand2_4 _30731_ (.A(_19919_),
    .B(_20117_),
    .Y(_08181_));
 sky130_fd_sc_hd__nand2_4 _30732_ (.A(_05366_),
    .B(_07232_),
    .Y(_08182_));
 sky130_fd_sc_hd__nor2_4 _30733_ (.A(_08181_),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__and2_1 _30734_ (.A(_08181_),
    .B(_08182_),
    .X(_08184_));
 sky130_fd_sc_hd__nand2_2 _30735_ (.A(_19936_),
    .B(\pcpi_mul.rs1[23] ),
    .Y(_08185_));
 sky130_fd_sc_hd__o21ai_2 _30736_ (.A1(_08183_),
    .A2(_08184_),
    .B1(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__or2_2 _30737_ (.A(_08181_),
    .B(_08182_),
    .X(_08187_));
 sky130_vsdinv _30738_ (.A(_08185_),
    .Y(_08188_));
 sky130_fd_sc_hd__nand2_4 _30739_ (.A(_08181_),
    .B(_08182_),
    .Y(_08189_));
 sky130_fd_sc_hd__nand3_4 _30740_ (.A(_08187_),
    .B(_08188_),
    .C(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand3_4 _30741_ (.A(_08180_),
    .B(_08186_),
    .C(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__o21ai_2 _30742_ (.A1(_08183_),
    .A2(_08184_),
    .B1(_08188_),
    .Y(_08192_));
 sky130_fd_sc_hd__nand3_2 _30743_ (.A(_08187_),
    .B(_08185_),
    .C(_08189_),
    .Y(_08193_));
 sky130_fd_sc_hd__a21oi_4 _30744_ (.A1(_08047_),
    .A2(_08043_),
    .B1(_08046_),
    .Y(_08194_));
 sky130_fd_sc_hd__nand3_4 _30745_ (.A(_08192_),
    .B(_08193_),
    .C(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__buf_4 _30746_ (.A(\pcpi_mul.rs1[21] ),
    .X(_08196_));
 sky130_fd_sc_hd__nand2_2 _30747_ (.A(_05235_),
    .B(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__a21o_1 _30748_ (.A1(_05477_),
    .A2(_20104_),
    .B1(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__nand2_2 _30749_ (.A(_19933_),
    .B(_08036_),
    .Y(_08199_));
 sky130_fd_sc_hd__a21o_1 _30750_ (.A1(_05387_),
    .A2(_08057_),
    .B1(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__nand2_2 _30751_ (.A(_05247_),
    .B(_08056_),
    .Y(_08201_));
 sky130_fd_sc_hd__a21oi_4 _30752_ (.A1(_08198_),
    .A2(_08200_),
    .B1(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__and3_2 _30753_ (.A(_08198_),
    .B(_08200_),
    .C(_08201_),
    .X(_08203_));
 sky130_fd_sc_hd__nor2_8 _30754_ (.A(_08202_),
    .B(_08203_),
    .Y(_08204_));
 sky130_fd_sc_hd__a21o_4 _30755_ (.A1(_08191_),
    .A2(_08195_),
    .B1(_08204_),
    .X(_08205_));
 sky130_fd_sc_hd__nand3_4 _30756_ (.A(_08204_),
    .B(_08191_),
    .C(_08195_),
    .Y(_08206_));
 sky130_fd_sc_hd__o21ai_4 _30757_ (.A1(_08064_),
    .A2(_08050_),
    .B1(_08068_),
    .Y(_08207_));
 sky130_fd_sc_hd__a21oi_1 _30758_ (.A1(_08205_),
    .A2(_08206_),
    .B1(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__and3_1 _30759_ (.A(_08186_),
    .B(_08180_),
    .C(_08190_),
    .X(_08209_));
 sky130_fd_sc_hd__nand2_1 _30760_ (.A(_08204_),
    .B(_08195_),
    .Y(_08210_));
 sky130_fd_sc_hd__o211a_4 _30761_ (.A1(_08209_),
    .A2(_08210_),
    .B1(_08207_),
    .C1(_08205_),
    .X(_08211_));
 sky130_fd_sc_hd__or2_1 _30762_ (.A(_08054_),
    .B(_08058_),
    .X(_08212_));
 sky130_fd_sc_hd__nand2_4 _30763_ (.A(_08062_),
    .B(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__o21ai_1 _30764_ (.A1(_08208_),
    .A2(_08211_),
    .B1(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__a21o_1 _30765_ (.A1(_08205_),
    .A2(_08206_),
    .B1(_08207_),
    .X(_08215_));
 sky130_vsdinv _30766_ (.A(_08213_),
    .Y(_08216_));
 sky130_fd_sc_hd__nand3_4 _30767_ (.A(_08205_),
    .B(_08207_),
    .C(_08206_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand3_1 _30768_ (.A(_08215_),
    .B(_08216_),
    .C(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__nand2_2 _30769_ (.A(_08214_),
    .B(_08218_),
    .Y(_08219_));
 sky130_fd_sc_hd__o21ai_2 _30770_ (.A1(_08175_),
    .A2(_08179_),
    .B1(_08219_),
    .Y(_08220_));
 sky130_fd_sc_hd__a22o_2 _30771_ (.A1(_08020_),
    .A2(_08139_),
    .B1(_08169_),
    .B2(_08174_),
    .X(_08221_));
 sky130_fd_sc_hd__nand2_2 _30772_ (.A(_08215_),
    .B(_08213_),
    .Y(_08222_));
 sky130_fd_sc_hd__o21ai_1 _30773_ (.A1(_08208_),
    .A2(_08211_),
    .B1(_08216_),
    .Y(_08223_));
 sky130_fd_sc_hd__o21ai_1 _30774_ (.A1(_08211_),
    .A2(_08222_),
    .B1(_08223_),
    .Y(_08224_));
 sky130_fd_sc_hd__o211ai_4 _30775_ (.A1(_08177_),
    .A2(_08178_),
    .B1(_08174_),
    .C1(_08169_),
    .Y(_08225_));
 sky130_fd_sc_hd__nand3_2 _30776_ (.A(_08221_),
    .B(_08224_),
    .C(_08225_),
    .Y(_08226_));
 sky130_fd_sc_hd__nand3_4 _30777_ (.A(_08220_),
    .B(_07959_),
    .C(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__a21oi_2 _30778_ (.A1(_08215_),
    .A2(_08217_),
    .B1(_08213_),
    .Y(_08228_));
 sky130_fd_sc_hd__nor2_2 _30779_ (.A(_08211_),
    .B(_08222_),
    .Y(_08229_));
 sky130_fd_sc_hd__o22ai_4 _30780_ (.A1(_08228_),
    .A2(_08229_),
    .B1(_08175_),
    .B2(_08179_),
    .Y(_08230_));
 sky130_fd_sc_hd__nand3_2 _30781_ (.A(_08221_),
    .B(_08225_),
    .C(_08219_),
    .Y(_08231_));
 sky130_vsdinv _30782_ (.A(_07959_),
    .Y(_08232_));
 sky130_fd_sc_hd__nand3_4 _30783_ (.A(_08230_),
    .B(_08231_),
    .C(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand2_1 _30784_ (.A(_08227_),
    .B(_08233_),
    .Y(_08234_));
 sky130_vsdinv _30785_ (.A(_08027_),
    .Y(_08235_));
 sky130_fd_sc_hd__a21o_1 _30786_ (.A1(_08080_),
    .A2(_08034_),
    .B1(_08235_),
    .X(_08236_));
 sky130_vsdinv _30787_ (.A(_08236_),
    .Y(_08237_));
 sky130_fd_sc_hd__nand2_4 _30788_ (.A(_08234_),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__nand3_2 _30789_ (.A(_08227_),
    .B(_08233_),
    .C(_08236_),
    .Y(_08239_));
 sky130_fd_sc_hd__buf_4 _30790_ (.A(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__nand2_1 _30791_ (.A(_08238_),
    .B(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__inv_8 _30792_ (.A(_05453_),
    .Y(_08242_));
 sky130_fd_sc_hd__buf_4 _30793_ (.A(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__a22oi_4 _30794_ (.A1(_19880_),
    .A2(_20158_),
    .B1(_06925_),
    .B2(_06472_),
    .Y(_08244_));
 sky130_fd_sc_hd__nand3_4 _30795_ (.A(_07087_),
    .B(_06636_),
    .C(_05664_),
    .Y(_08245_));
 sky130_fd_sc_hd__nor2_8 _30796_ (.A(_06247_),
    .B(_08245_),
    .Y(_08246_));
 sky130_fd_sc_hd__o22ai_4 _30797_ (.A1(_06528_),
    .A2(net442),
    .B1(_08244_),
    .B2(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__buf_6 _30798_ (.A(_07827_),
    .X(_08248_));
 sky130_fd_sc_hd__a22oi_4 _30799_ (.A1(_07482_),
    .A2(_05300_),
    .B1(_08248_),
    .B2(_20168_),
    .Y(_08249_));
 sky130_fd_sc_hd__o21ai_4 _30800_ (.A1(_07978_),
    .A2(_08249_),
    .B1(_07974_),
    .Y(_08250_));
 sky130_fd_sc_hd__nand2_2 _30801_ (.A(_07893_),
    .B(_20151_),
    .Y(_08251_));
 sky130_vsdinv _30802_ (.A(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__a22o_2 _30803_ (.A1(_07446_),
    .A2(_07417_),
    .B1(_19886_),
    .B2(_05696_),
    .X(_08253_));
 sky130_fd_sc_hd__o211ai_2 _30804_ (.A1(_06248_),
    .A2(_08245_),
    .B1(_08252_),
    .C1(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__nand3_4 _30805_ (.A(_08247_),
    .B(_08250_),
    .C(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__o21ai_4 _30806_ (.A1(_08244_),
    .A2(_08246_),
    .B1(_08252_),
    .Y(_08256_));
 sky130_fd_sc_hd__o21ai_2 _30807_ (.A1(_07972_),
    .A2(_07975_),
    .B1(_07978_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand2_4 _30808_ (.A(_08257_),
    .B(_07976_),
    .Y(_08258_));
 sky130_fd_sc_hd__o211ai_4 _30809_ (.A1(_06248_),
    .A2(_08245_),
    .B1(_08251_),
    .C1(_08253_),
    .Y(_08259_));
 sky130_fd_sc_hd__nand3_4 _30810_ (.A(_08256_),
    .B(_08258_),
    .C(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__nor2_2 _30811_ (.A(_07898_),
    .B(_07892_),
    .Y(_08261_));
 sky130_fd_sc_hd__o2bb2ai_4 _30812_ (.A1_N(_08255_),
    .A2_N(_08260_),
    .B1(_07891_),
    .B2(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__a21oi_4 _30813_ (.A1(_07899_),
    .A2(_07898_),
    .B1(_07892_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand3b_4 _30814_ (.A_N(_08263_),
    .B(_08260_),
    .C(_08255_),
    .Y(_08264_));
 sky130_fd_sc_hd__nand2_2 _30815_ (.A(_07919_),
    .B(_07905_),
    .Y(_08265_));
 sky130_fd_sc_hd__a21oi_4 _30816_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__o211a_4 _30817_ (.A1(_07918_),
    .A2(_07914_),
    .B1(_08264_),
    .C1(_08262_),
    .X(_08267_));
 sky130_fd_sc_hd__a22oi_4 _30818_ (.A1(_07102_),
    .A2(_05555_),
    .B1(_06545_),
    .B2(_05822_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_2 _30819_ (.A(\pcpi_mul.rs2[14] ),
    .B(_05554_),
    .Y(_08269_));
 sky130_fd_sc_hd__nand2_2 _30820_ (.A(_06606_),
    .B(_05670_),
    .Y(_08270_));
 sky130_fd_sc_hd__nor2_4 _30821_ (.A(_08269_),
    .B(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__nand2_2 _30822_ (.A(_07785_),
    .B(_06153_),
    .Y(_08272_));
 sky130_fd_sc_hd__o21bai_4 _30823_ (.A1(_08268_),
    .A2(_08271_),
    .B1_N(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__nand3b_4 _30824_ (.A_N(_08269_),
    .B(_06207_),
    .C(_06841_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand2_2 _30825_ (.A(_08269_),
    .B(_08270_),
    .Y(_08275_));
 sky130_fd_sc_hd__nand3_4 _30826_ (.A(_08274_),
    .B(_08275_),
    .C(_08272_),
    .Y(_08276_));
 sky130_fd_sc_hd__nor2_2 _30827_ (.A(_07927_),
    .B(_07923_),
    .Y(_08277_));
 sky130_fd_sc_hd__o2bb2ai_4 _30828_ (.A1_N(_08273_),
    .A2_N(_08276_),
    .B1(_07926_),
    .B2(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__a21oi_2 _30829_ (.A1(_07928_),
    .A2(_07931_),
    .B1(_07926_),
    .Y(_08279_));
 sky130_fd_sc_hd__nand3_4 _30830_ (.A(_08273_),
    .B(_08276_),
    .C(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__nand2_1 _30831_ (.A(_08278_),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__a22oi_4 _30832_ (.A1(_19901_),
    .A2(_06309_),
    .B1(_19905_),
    .B2(_07661_),
    .Y(_08282_));
 sky130_fd_sc_hd__nand2_1 _30833_ (.A(_06622_),
    .B(_20137_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_1 _30834_ (.A(_05656_),
    .B(_06142_),
    .Y(_08284_));
 sky130_fd_sc_hd__nor2_1 _30835_ (.A(_08283_),
    .B(_08284_),
    .Y(_08285_));
 sky130_fd_sc_hd__nand2_2 _30836_ (.A(_19908_),
    .B(_06294_),
    .Y(_08286_));
 sky130_fd_sc_hd__o21bai_2 _30837_ (.A1(_08282_),
    .A2(_08285_),
    .B1_N(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__nand3b_2 _30838_ (.A_N(_08283_),
    .B(_06631_),
    .C(_07503_),
    .Y(_08288_));
 sky130_fd_sc_hd__nand2_1 _30839_ (.A(_08283_),
    .B(_08284_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand3_2 _30840_ (.A(_08288_),
    .B(_08289_),
    .C(_08286_),
    .Y(_08290_));
 sky130_fd_sc_hd__nand2_4 _30841_ (.A(_08287_),
    .B(_08290_),
    .Y(_08291_));
 sky130_vsdinv _30842_ (.A(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand2_1 _30843_ (.A(_08281_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__nand3_1 _30844_ (.A(_08278_),
    .B(_08280_),
    .C(_08291_),
    .Y(_08294_));
 sky130_fd_sc_hd__nand2_2 _30845_ (.A(_08293_),
    .B(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__o21ai_2 _30846_ (.A1(_08266_),
    .A2(_08267_),
    .B1(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__a21o_1 _30847_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08265_),
    .X(_08297_));
 sky130_fd_sc_hd__nand2_1 _30848_ (.A(_08281_),
    .B(_08291_),
    .Y(_08298_));
 sky130_fd_sc_hd__nand3_2 _30849_ (.A(_08292_),
    .B(_08280_),
    .C(_08278_),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_4 _30850_ (.A(_08298_),
    .B(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__nand3_4 _30851_ (.A(_08265_),
    .B(_08262_),
    .C(_08264_),
    .Y(_08301_));
 sky130_fd_sc_hd__nand3_4 _30852_ (.A(_08297_),
    .B(_08300_),
    .C(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__nand3_4 _30853_ (.A(_08296_),
    .B(_07985_),
    .C(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__nor2_2 _30854_ (.A(_08291_),
    .B(_08281_),
    .Y(_08304_));
 sky130_fd_sc_hd__a21oi_2 _30855_ (.A1(_08278_),
    .A2(_08280_),
    .B1(_08292_),
    .Y(_08305_));
 sky130_fd_sc_hd__o22ai_4 _30856_ (.A1(_08304_),
    .A2(_08305_),
    .B1(_08266_),
    .B2(_08267_),
    .Y(_08306_));
 sky130_fd_sc_hd__nand3_4 _30857_ (.A(_08297_),
    .B(_08295_),
    .C(_08301_),
    .Y(_08307_));
 sky130_fd_sc_hd__nand3_4 _30858_ (.A(_08306_),
    .B(_07984_),
    .C(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__nand2_1 _30859_ (.A(_08303_),
    .B(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__o21ai_4 _30860_ (.A1(_07950_),
    .A2(_07917_),
    .B1(_07954_),
    .Y(_08310_));
 sky130_vsdinv _30861_ (.A(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__nand2_2 _30862_ (.A(_08309_),
    .B(_08311_),
    .Y(_08312_));
 sky130_fd_sc_hd__nand3_2 _30863_ (.A(_08303_),
    .B(_08308_),
    .C(_08310_),
    .Y(_08313_));
 sky130_fd_sc_hd__nand2_2 _30864_ (.A(_19862_),
    .B(_05145_),
    .Y(_08314_));
 sky130_fd_sc_hd__clkbuf_4 _30865_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08315_));
 sky130_fd_sc_hd__nand2_2 _30866_ (.A(_08315_),
    .B(_20176_),
    .Y(_08316_));
 sky130_fd_sc_hd__nor2_4 _30867_ (.A(_08314_),
    .B(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__and2_1 _30868_ (.A(_08314_),
    .B(_08316_),
    .X(_08318_));
 sky130_fd_sc_hd__nor2_4 _30869_ (.A(_07822_),
    .B(_05126_),
    .Y(_08319_));
 sky130_fd_sc_hd__o21bai_2 _30870_ (.A1(_08317_),
    .A2(_08318_),
    .B1_N(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__nand2_2 _30871_ (.A(_08314_),
    .B(_08316_),
    .Y(_08321_));
 sky130_fd_sc_hd__nand3b_4 _30872_ (.A_N(_08317_),
    .B(_08319_),
    .C(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__a21o_4 _30873_ (.A1(_08320_),
    .A2(_08322_),
    .B1(_07970_),
    .X(_08323_));
 sky130_fd_sc_hd__nand3_4 _30874_ (.A(_08320_),
    .B(_08322_),
    .C(_07970_),
    .Y(_08324_));
 sky130_fd_sc_hd__nand2_2 _30875_ (.A(_08323_),
    .B(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__buf_6 _30876_ (.A(_07481_),
    .X(_08326_));
 sky130_fd_sc_hd__a22oi_4 _30877_ (.A1(_08326_),
    .A2(_05182_),
    .B1(_07354_),
    .B2(_05283_),
    .Y(_08327_));
 sky130_fd_sc_hd__nand3_4 _30878_ (.A(_07482_),
    .B(_07354_),
    .C(_20168_),
    .Y(_08328_));
 sky130_fd_sc_hd__nor2_1 _30879_ (.A(_05253_),
    .B(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__a211o_1 _30880_ (.A1(_19878_),
    .A2(_20163_),
    .B1(_08327_),
    .C1(_08329_),
    .X(_08330_));
 sky130_fd_sc_hd__nand2_2 _30881_ (.A(_19877_),
    .B(_05286_),
    .Y(_08331_));
 sky130_fd_sc_hd__o21bai_2 _30882_ (.A1(_08327_),
    .A2(_08329_),
    .B1_N(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand2_4 _30883_ (.A(_08330_),
    .B(_08332_),
    .Y(_08333_));
 sky130_vsdinv _30884_ (.A(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__nand2_2 _30885_ (.A(_08325_),
    .B(_08334_),
    .Y(_08335_));
 sky130_fd_sc_hd__nand3_4 _30886_ (.A(_08323_),
    .B(_08324_),
    .C(_08333_),
    .Y(_08336_));
 sky130_fd_sc_hd__a21boi_1 _30887_ (.A1(_08335_),
    .A2(_08336_),
    .B1_N(_07982_),
    .Y(_08337_));
 sky130_fd_sc_hd__a31o_1 _30888_ (.A1(_08323_),
    .A2(_08324_),
    .A3(_08333_),
    .B1(_07982_),
    .X(_08338_));
 sky130_fd_sc_hd__a21oi_4 _30889_ (.A1(_08325_),
    .A2(_08334_),
    .B1(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__or2_4 _30890_ (.A(_08337_),
    .B(_08339_),
    .X(_08340_));
 sky130_vsdinv _30891_ (.A(_08340_),
    .Y(_08341_));
 sky130_fd_sc_hd__a21oi_2 _30892_ (.A1(_08312_),
    .A2(_08313_),
    .B1(_08341_),
    .Y(_08342_));
 sky130_fd_sc_hd__a21oi_4 _30893_ (.A1(_08303_),
    .A2(_08308_),
    .B1(_08310_),
    .Y(_08343_));
 sky130_fd_sc_hd__and3_2 _30894_ (.A(_08303_),
    .B(_08308_),
    .C(_08310_),
    .X(_08344_));
 sky130_fd_sc_hd__nor3_4 _30895_ (.A(_08340_),
    .B(_08343_),
    .C(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__o22ai_4 _30896_ (.A1(_08098_),
    .A2(_08097_),
    .B1(_08342_),
    .B2(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__o21ai_2 _30897_ (.A1(_08343_),
    .A2(_08344_),
    .B1(_08340_),
    .Y(_08347_));
 sky130_vsdinv _30898_ (.A(_07988_),
    .Y(_08348_));
 sky130_fd_sc_hd__nand3_2 _30899_ (.A(_08312_),
    .B(_08341_),
    .C(_08313_),
    .Y(_08349_));
 sky130_fd_sc_hd__nand3_4 _30900_ (.A(_08347_),
    .B(_08348_),
    .C(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__nand3_2 _30901_ (.A(_08241_),
    .B(_08346_),
    .C(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__nand2_1 _30902_ (.A(_08346_),
    .B(_08350_),
    .Y(_08352_));
 sky130_fd_sc_hd__nand3_2 _30903_ (.A(_08352_),
    .B(_08238_),
    .C(_08240_),
    .Y(_08353_));
 sky130_fd_sc_hd__a31oi_4 _30904_ (.A1(_08096_),
    .A2(_08106_),
    .A3(_08101_),
    .B1(_07991_),
    .Y(_08354_));
 sky130_fd_sc_hd__nand3_4 _30905_ (.A(_08351_),
    .B(_08353_),
    .C(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__a21oi_1 _30906_ (.A1(_08227_),
    .A2(_08233_),
    .B1(_08236_),
    .Y(_08356_));
 sky130_fd_sc_hd__and3_1 _30907_ (.A(_08227_),
    .B(_08233_),
    .C(_08236_),
    .X(_08357_));
 sky130_fd_sc_hd__o2bb2ai_2 _30908_ (.A1_N(_08346_),
    .A2_N(_08350_),
    .B1(_08356_),
    .B2(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__o21bai_2 _30909_ (.A1(_08092_),
    .A2(_08108_),
    .B1_N(_07991_),
    .Y(_08359_));
 sky130_fd_sc_hd__nand2_1 _30910_ (.A(_08347_),
    .B(_08348_),
    .Y(_08360_));
 sky130_fd_sc_hd__o2111ai_4 _30911_ (.A1(_08345_),
    .A2(_08360_),
    .B1(_08240_),
    .C1(_08346_),
    .D1(_08238_),
    .Y(_08361_));
 sky130_fd_sc_hd__nand3_4 _30912_ (.A(_08358_),
    .B(_08359_),
    .C(_08361_),
    .Y(_08362_));
 sky130_vsdinv _30913_ (.A(_08077_),
    .Y(_08363_));
 sky130_fd_sc_hd__nand2_4 _30914_ (.A(_08363_),
    .B(_08072_),
    .Y(_08364_));
 sky130_fd_sc_hd__nand2_4 _30915_ (.A(_08101_),
    .B(_08089_),
    .Y(_08365_));
 sky130_fd_sc_hd__xor2_4 _30916_ (.A(_08364_),
    .B(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__a21o_1 _30917_ (.A1(_08355_),
    .A2(_08362_),
    .B1(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__nand3_4 _30918_ (.A(_08355_),
    .B(_08362_),
    .C(_08366_),
    .Y(_08368_));
 sky130_vsdinv _30919_ (.A(_08113_),
    .Y(_08369_));
 sky130_fd_sc_hd__o21ai_2 _30920_ (.A1(_08105_),
    .A2(_08369_),
    .B1(_08112_),
    .Y(_08370_));
 sky130_fd_sc_hd__nand3_4 _30921_ (.A(_08367_),
    .B(_08368_),
    .C(_08370_),
    .Y(_08371_));
 sky130_vsdinv _30922_ (.A(_08365_),
    .Y(_08372_));
 sky130_fd_sc_hd__nor2_1 _30923_ (.A(_08364_),
    .B(_08372_),
    .Y(_08373_));
 sky130_vsdinv _30924_ (.A(_08364_),
    .Y(_08374_));
 sky130_fd_sc_hd__nor2_1 _30925_ (.A(_08374_),
    .B(_08365_),
    .Y(_08375_));
 sky130_fd_sc_hd__o2bb2ai_2 _30926_ (.A1_N(_08362_),
    .A2_N(_08355_),
    .B1(_08373_),
    .B2(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__a21oi_4 _30927_ (.A1(_08111_),
    .A2(_08113_),
    .B1(_08109_),
    .Y(_08377_));
 sky130_fd_sc_hd__nand2_1 _30928_ (.A(_08372_),
    .B(_08374_),
    .Y(_08378_));
 sky130_fd_sc_hd__nand2_2 _30929_ (.A(_08365_),
    .B(_08364_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand2_2 _30930_ (.A(_08378_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__nand3_4 _30931_ (.A(_08355_),
    .B(_08380_),
    .C(_08362_),
    .Y(_08381_));
 sky130_fd_sc_hd__nand3_4 _30932_ (.A(_08376_),
    .B(_08377_),
    .C(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__buf_2 _30933_ (.A(_07889_),
    .X(_08383_));
 sky130_fd_sc_hd__a21oi_2 _30934_ (.A1(_08371_),
    .A2(_08382_),
    .B1(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand3_1 _30935_ (.A(_08371_),
    .B(_08382_),
    .C(_08383_),
    .Y(_08385_));
 sky130_fd_sc_hd__nand2_1 _30936_ (.A(_08125_),
    .B(_07865_),
    .Y(_08386_));
 sky130_fd_sc_hd__nand3_2 _30937_ (.A(_08385_),
    .B(_08124_),
    .C(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__nand2_1 _30938_ (.A(_08371_),
    .B(_08382_),
    .Y(_08388_));
 sky130_fd_sc_hd__nand2_1 _30939_ (.A(_08388_),
    .B(_08383_),
    .Y(_08389_));
 sky130_fd_sc_hd__nand2_1 _30940_ (.A(_08386_),
    .B(_08124_),
    .Y(_08390_));
 sky130_fd_sc_hd__nand3b_2 _30941_ (.A_N(_08383_),
    .B(_08371_),
    .C(_08382_),
    .Y(_08391_));
 sky130_fd_sc_hd__nand3_2 _30942_ (.A(_08389_),
    .B(_08390_),
    .C(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__o21a_1 _30943_ (.A1(_08384_),
    .A2(_08387_),
    .B1(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__a21oi_1 _30944_ (.A1(_08138_),
    .A2(_08132_),
    .B1(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__and3_1 _30945_ (.A(_08138_),
    .B(_08132_),
    .C(_08393_),
    .X(_08395_));
 sky130_fd_sc_hd__or2_1 _30946_ (.A(_08394_),
    .B(_08395_),
    .X(_02642_));
 sky130_fd_sc_hd__nand3_4 _30947_ (.A(_08238_),
    .B(_08346_),
    .C(_08240_),
    .Y(_08396_));
 sky130_fd_sc_hd__nand2_1 _30948_ (.A(_08396_),
    .B(_08350_),
    .Y(_08397_));
 sky130_fd_sc_hd__a22oi_4 _30949_ (.A1(_07660_),
    .A2(_06816_),
    .B1(_05413_),
    .B2(_06979_),
    .Y(_08398_));
 sky130_fd_sc_hd__nor2_4 _30950_ (.A(_08039_),
    .B(_08149_),
    .Y(_08399_));
 sky130_fd_sc_hd__nand2_2 _30951_ (.A(_05865_),
    .B(_07249_),
    .Y(_08400_));
 sky130_fd_sc_hd__o21ai_2 _30952_ (.A1(_08398_),
    .A2(_08399_),
    .B1(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__o21ai_2 _30953_ (.A1(_08286_),
    .A2(_08282_),
    .B1(_08288_),
    .Y(_08402_));
 sky130_vsdinv _30954_ (.A(_08400_),
    .Y(_08403_));
 sky130_fd_sc_hd__a22o_2 _30955_ (.A1(_06478_),
    .A2(_06816_),
    .B1(_06097_),
    .B2(_07251_),
    .X(_08404_));
 sky130_fd_sc_hd__o211ai_4 _30956_ (.A1(_08040_),
    .A2(_08149_),
    .B1(_08403_),
    .C1(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__nand3_4 _30957_ (.A(_08401_),
    .B(_08402_),
    .C(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__o21ai_2 _30958_ (.A1(_08398_),
    .A2(_08399_),
    .B1(_08403_),
    .Y(_08407_));
 sky130_fd_sc_hd__o21ai_1 _30959_ (.A1(_08283_),
    .A2(_08284_),
    .B1(_08286_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand2_1 _30960_ (.A(_08408_),
    .B(_08289_),
    .Y(_08409_));
 sky130_fd_sc_hd__o211ai_4 _30961_ (.A1(_08040_),
    .A2(_08149_),
    .B1(_08400_),
    .C1(_08404_),
    .Y(_08410_));
 sky130_fd_sc_hd__nand3_4 _30962_ (.A(_08407_),
    .B(_08409_),
    .C(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__nor2_4 _30963_ (.A(_08150_),
    .B(_08145_),
    .Y(_08412_));
 sky130_fd_sc_hd__o2bb2ai_4 _30964_ (.A1_N(_08406_),
    .A2_N(_08411_),
    .B1(_08143_),
    .B2(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__nor2_2 _30965_ (.A(_08143_),
    .B(_08412_),
    .Y(_08414_));
 sky130_fd_sc_hd__nand3_4 _30966_ (.A(_08406_),
    .B(_08411_),
    .C(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2_1 _30967_ (.A(_08280_),
    .B(_08291_),
    .Y(_08416_));
 sky130_fd_sc_hd__nand2_4 _30968_ (.A(_08416_),
    .B(_08278_),
    .Y(_08417_));
 sky130_fd_sc_hd__a21oi_4 _30969_ (.A1(_08413_),
    .A2(_08415_),
    .B1(_08417_),
    .Y(_08418_));
 sky130_fd_sc_hd__nand2_1 _30970_ (.A(_08411_),
    .B(_08414_),
    .Y(_08419_));
 sky130_vsdinv _30971_ (.A(_08406_),
    .Y(_08420_));
 sky130_fd_sc_hd__o211a_1 _30972_ (.A1(_08419_),
    .A2(_08420_),
    .B1(_08413_),
    .C1(_08417_),
    .X(_08421_));
 sky130_fd_sc_hd__and2_2 _30973_ (.A(_08167_),
    .B(_08154_),
    .X(_08422_));
 sky130_fd_sc_hd__o21ai_4 _30974_ (.A1(_08418_),
    .A2(_08421_),
    .B1(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__a21o_1 _30975_ (.A1(_08413_),
    .A2(_08415_),
    .B1(_08417_),
    .X(_08424_));
 sky130_fd_sc_hd__nand3_4 _30976_ (.A(_08417_),
    .B(_08413_),
    .C(_08415_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand3b_4 _30977_ (.A_N(_08422_),
    .B(_08424_),
    .C(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand2_1 _30978_ (.A(_08173_),
    .B(_08171_),
    .Y(_08427_));
 sky130_fd_sc_hd__nand2_1 _30979_ (.A(_08427_),
    .B(_08172_),
    .Y(_08428_));
 sky130_fd_sc_hd__a21boi_4 _30980_ (.A1(_08423_),
    .A2(_08426_),
    .B1_N(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__nor2_1 _30981_ (.A(_08171_),
    .B(_08165_),
    .Y(_08430_));
 sky130_fd_sc_hd__o211a_2 _30982_ (.A1(_08168_),
    .A2(_08430_),
    .B1(_08426_),
    .C1(_08423_),
    .X(_08431_));
 sky130_fd_sc_hd__and4_2 _30983_ (.A(_05302_),
    .B(_05366_),
    .C(_07722_),
    .D(_20113_),
    .X(_08432_));
 sky130_fd_sc_hd__clkbuf_4 _30984_ (.A(_07232_),
    .X(_08433_));
 sky130_fd_sc_hd__a22o_2 _30985_ (.A1(_05228_),
    .A2(_08433_),
    .B1(_05312_),
    .B2(_07548_),
    .X(_08434_));
 sky130_vsdinv _30986_ (.A(\pcpi_mul.rs1[24] ),
    .Y(_08435_));
 sky130_fd_sc_hd__nor2_4 _30987_ (.A(_04836_),
    .B(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__nand3b_4 _30988_ (.A_N(_08432_),
    .B(_08434_),
    .C(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__a22oi_4 _30989_ (.A1(_05213_),
    .A2(_07233_),
    .B1(_05298_),
    .B2(_08053_),
    .Y(_08438_));
 sky130_fd_sc_hd__o21bai_4 _30990_ (.A1(_08438_),
    .A2(_08432_),
    .B1_N(_08436_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand2_1 _30991_ (.A(_08437_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_4 _30992_ (.A1(_08188_),
    .A2(_08189_),
    .B1(_08183_),
    .Y(_08441_));
 sky130_fd_sc_hd__nand2_4 _30993_ (.A(_08440_),
    .B(_08441_),
    .Y(_08442_));
 sky130_vsdinv _30994_ (.A(_08441_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand3_4 _30995_ (.A(_08443_),
    .B(_08437_),
    .C(_08439_),
    .Y(_08444_));
 sky130_fd_sc_hd__buf_2 _30996_ (.A(\pcpi_mul.rs1[23] ),
    .X(_08445_));
 sky130_fd_sc_hd__clkbuf_4 _30997_ (.A(_08445_),
    .X(_08446_));
 sky130_fd_sc_hd__buf_4 _30998_ (.A(\pcpi_mul.rs1[22] ),
    .X(_08447_));
 sky130_fd_sc_hd__nand2_2 _30999_ (.A(_05173_),
    .B(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__a21o_2 _31000_ (.A1(_19934_),
    .A2(_08446_),
    .B1(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__clkbuf_4 _31001_ (.A(_08036_),
    .X(_08450_));
 sky130_fd_sc_hd__nand2_2 _31002_ (.A(_05570_),
    .B(_08445_),
    .Y(_08451_));
 sky130_fd_sc_hd__a21o_2 _31003_ (.A1(_05240_),
    .A2(_08450_),
    .B1(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__buf_6 _31004_ (.A(_08196_),
    .X(_08453_));
 sky130_fd_sc_hd__nand2_4 _31005_ (.A(_05692_),
    .B(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand3_4 _31006_ (.A(_08449_),
    .B(_08452_),
    .C(_08454_),
    .Y(_08455_));
 sky130_vsdinv _31007_ (.A(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__a21oi_4 _31008_ (.A1(_08449_),
    .A2(_08452_),
    .B1(_08454_),
    .Y(_08457_));
 sky130_fd_sc_hd__o2bb2ai_2 _31009_ (.A1_N(_08442_),
    .A2_N(_08444_),
    .B1(_08456_),
    .B2(_08457_),
    .Y(_08458_));
 sky130_vsdinv _31010_ (.A(_08186_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand2_1 _31011_ (.A(_08180_),
    .B(_08190_),
    .Y(_08460_));
 sky130_fd_sc_hd__o2bb2ai_2 _31012_ (.A1_N(_08204_),
    .A2_N(_08195_),
    .B1(_08459_),
    .B2(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__nor2_2 _31013_ (.A(_08457_),
    .B(_08456_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand3_2 _31014_ (.A(_08462_),
    .B(_08442_),
    .C(_08444_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand3_4 _31015_ (.A(_08458_),
    .B(_08461_),
    .C(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__nand2_1 _31016_ (.A(_08442_),
    .B(_08444_),
    .Y(_08465_));
 sky130_fd_sc_hd__nand2_2 _31017_ (.A(_08465_),
    .B(_08462_),
    .Y(_08466_));
 sky130_fd_sc_hd__a21oi_4 _31018_ (.A1(_08204_),
    .A2(_08195_),
    .B1(_08209_),
    .Y(_08467_));
 sky130_fd_sc_hd__a21o_1 _31019_ (.A1(_08449_),
    .A2(_08452_),
    .B1(_08454_),
    .X(_08468_));
 sky130_fd_sc_hd__nand2_4 _31020_ (.A(_08468_),
    .B(_08455_),
    .Y(_08469_));
 sky130_fd_sc_hd__nand3_4 _31021_ (.A(_08442_),
    .B(_08444_),
    .C(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__nor2_4 _31022_ (.A(_08197_),
    .B(_08199_),
    .Y(_08471_));
 sky130_fd_sc_hd__nor2_8 _31023_ (.A(_08471_),
    .B(_08202_),
    .Y(_08472_));
 sky130_fd_sc_hd__a31oi_4 _31024_ (.A1(_08466_),
    .A2(_08467_),
    .A3(_08470_),
    .B1(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__nand3_4 _31025_ (.A(_08466_),
    .B(_08467_),
    .C(_08470_),
    .Y(_08474_));
 sky130_fd_sc_hd__a21boi_4 _31026_ (.A1(_08474_),
    .A2(_08464_),
    .B1_N(_08472_),
    .Y(_08475_));
 sky130_fd_sc_hd__a21oi_4 _31027_ (.A1(_08464_),
    .A2(_08473_),
    .B1(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__o21ai_2 _31028_ (.A1(_08429_),
    .A2(_08431_),
    .B1(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__a21boi_2 _31029_ (.A1(_08308_),
    .A2(_08310_),
    .B1_N(_08303_),
    .Y(_08478_));
 sky130_fd_sc_hd__a22o_1 _31030_ (.A1(_08172_),
    .A2(_08427_),
    .B1(_08423_),
    .B2(_08426_),
    .X(_08479_));
 sky130_fd_sc_hd__nand2_1 _31031_ (.A(_08474_),
    .B(_08464_),
    .Y(_08480_));
 sky130_fd_sc_hd__nand2_1 _31032_ (.A(_08480_),
    .B(_08472_),
    .Y(_08481_));
 sky130_fd_sc_hd__nand2_1 _31033_ (.A(_08473_),
    .B(_08464_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand2_1 _31034_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__nand3b_4 _31035_ (.A_N(_08428_),
    .B(_08426_),
    .C(_08423_),
    .Y(_08484_));
 sky130_fd_sc_hd__nand3_2 _31036_ (.A(_08479_),
    .B(_08483_),
    .C(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nand3_4 _31037_ (.A(_08477_),
    .B(_08478_),
    .C(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__nor2_2 _31038_ (.A(_08472_),
    .B(_08480_),
    .Y(_08487_));
 sky130_fd_sc_hd__o22ai_4 _31039_ (.A1(_08487_),
    .A2(_08475_),
    .B1(_08429_),
    .B2(_08431_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand3_2 _31040_ (.A(_08479_),
    .B(_08476_),
    .C(_08484_),
    .Y(_08489_));
 sky130_fd_sc_hd__nand2_1 _31041_ (.A(_08308_),
    .B(_08310_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_1 _31042_ (.A(_08490_),
    .B(_08303_),
    .Y(_08491_));
 sky130_fd_sc_hd__nand3_4 _31043_ (.A(_08488_),
    .B(_08489_),
    .C(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__nand2_4 _31044_ (.A(_08486_),
    .B(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__a21oi_4 _31045_ (.A1(_08221_),
    .A2(_08219_),
    .B1(_08179_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_8 _31046_ (.A(_08493_),
    .B(_08494_),
    .Y(_08495_));
 sky130_vsdinv _31047_ (.A(_08494_),
    .Y(_08496_));
 sky130_fd_sc_hd__nand3_4 _31048_ (.A(_08496_),
    .B(_08486_),
    .C(_08492_),
    .Y(_08497_));
 sky130_fd_sc_hd__clkbuf_4 _31049_ (.A(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__nand2_1 _31050_ (.A(_08255_),
    .B(_08263_),
    .Y(_08499_));
 sky130_fd_sc_hd__a22oi_4 _31051_ (.A1(_07289_),
    .A2(_20156_),
    .B1(_07449_),
    .B2(_05463_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand3_4 _31052_ (.A(_19880_),
    .B(_06925_),
    .C(_06472_),
    .Y(_08501_));
 sky130_fd_sc_hd__nor2_8 _31053_ (.A(_08242_),
    .B(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__nand2_2 _31054_ (.A(_07893_),
    .B(_05689_),
    .Y(_08503_));
 sky130_fd_sc_hd__o21ai_2 _31055_ (.A1(_08500_),
    .A2(_08502_),
    .B1(_08503_),
    .Y(_08504_));
 sky130_vsdinv _31056_ (.A(_08503_),
    .Y(_08505_));
 sky130_fd_sc_hd__a22o_4 _31057_ (.A1(_07289_),
    .A2(_20156_),
    .B1(_07291_),
    .B2(_05463_),
    .X(_08506_));
 sky130_fd_sc_hd__o211ai_4 _31058_ (.A1(net442),
    .A2(_08501_),
    .B1(_08505_),
    .C1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__o22ai_4 _31059_ (.A1(_05253_),
    .A2(_08328_),
    .B1(_08331_),
    .B2(_08327_),
    .Y(_08508_));
 sky130_fd_sc_hd__nand3_4 _31060_ (.A(_08504_),
    .B(_08507_),
    .C(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__o21ai_2 _31061_ (.A1(_08500_),
    .A2(_08502_),
    .B1(_08505_),
    .Y(_08510_));
 sky130_fd_sc_hd__o22a_2 _31062_ (.A1(_05253_),
    .A2(_08328_),
    .B1(_08331_),
    .B2(_08327_),
    .X(_08511_));
 sky130_fd_sc_hd__o211ai_4 _31063_ (.A1(net442),
    .A2(_08501_),
    .B1(_08503_),
    .C1(_08506_),
    .Y(_08512_));
 sky130_fd_sc_hd__nand3_4 _31064_ (.A(_08510_),
    .B(_08511_),
    .C(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__nor2_4 _31065_ (.A(_08252_),
    .B(_08246_),
    .Y(_08514_));
 sky130_fd_sc_hd__o2bb2ai_4 _31066_ (.A1_N(_08509_),
    .A2_N(_08513_),
    .B1(_08244_),
    .B2(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__nor2_4 _31067_ (.A(_08244_),
    .B(_08514_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand3_4 _31068_ (.A(_08513_),
    .B(_08509_),
    .C(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__a22oi_4 _31069_ (.A1(_08260_),
    .A2(_08499_),
    .B1(_08515_),
    .B2(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__a31oi_4 _31070_ (.A1(_08256_),
    .A2(_08258_),
    .A3(_08259_),
    .B1(_08263_),
    .Y(_08519_));
 sky130_vsdinv _31071_ (.A(_08255_),
    .Y(_08520_));
 sky130_fd_sc_hd__o211a_1 _31072_ (.A1(_08519_),
    .A2(_08520_),
    .B1(_08517_),
    .C1(_08515_),
    .X(_08521_));
 sky130_fd_sc_hd__nand2_4 _31073_ (.A(_19892_),
    .B(_05670_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand2_4 _31074_ (.A(_06606_),
    .B(_05998_),
    .Y(_08523_));
 sky130_fd_sc_hd__nor2_8 _31075_ (.A(_08522_),
    .B(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__nand2_2 _31076_ (.A(\pcpi_mul.rs2[12] ),
    .B(_20137_),
    .Y(_08525_));
 sky130_vsdinv _31077_ (.A(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_2 _31078_ (.A(_08522_),
    .B(_08523_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_2 _31079_ (.A(_08526_),
    .B(_08527_),
    .Y(_08528_));
 sky130_fd_sc_hd__o21ai_2 _31080_ (.A1(_08272_),
    .A2(_08268_),
    .B1(_08274_),
    .Y(_08529_));
 sky130_fd_sc_hd__buf_8 _31081_ (.A(_06153_),
    .X(_08530_));
 sky130_fd_sc_hd__a22oi_4 _31082_ (.A1(_06544_),
    .A2(_20146_),
    .B1(_06546_),
    .B2(_08530_),
    .Y(_08531_));
 sky130_fd_sc_hd__o21ai_2 _31083_ (.A1(_08531_),
    .A2(_08524_),
    .B1(_08525_),
    .Y(_08532_));
 sky130_fd_sc_hd__o211ai_4 _31084_ (.A1(_08524_),
    .A2(_08528_),
    .B1(_08529_),
    .C1(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__o21ai_2 _31085_ (.A1(_08531_),
    .A2(_08524_),
    .B1(_08526_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand3b_4 _31086_ (.A_N(_08522_),
    .B(_06546_),
    .C(_08530_),
    .Y(_08535_));
 sky130_fd_sc_hd__nand3_2 _31087_ (.A(_08535_),
    .B(_08527_),
    .C(_08525_),
    .Y(_08536_));
 sky130_vsdinv _31088_ (.A(_08272_),
    .Y(_08537_));
 sky130_fd_sc_hd__a21oi_2 _31089_ (.A1(_08537_),
    .A2(_08275_),
    .B1(_08271_),
    .Y(_08538_));
 sky130_fd_sc_hd__nand3_4 _31090_ (.A(_08534_),
    .B(_08536_),
    .C(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__a22oi_4 _31091_ (.A1(_06118_),
    .A2(_20135_),
    .B1(_06045_),
    .B2(_06718_),
    .Y(_08540_));
 sky130_fd_sc_hd__nand2_2 _31092_ (.A(_06117_),
    .B(_06142_),
    .Y(_08541_));
 sky130_fd_sc_hd__nand2_1 _31093_ (.A(_06106_),
    .B(_06294_),
    .Y(_08542_));
 sky130_fd_sc_hd__nor2_1 _31094_ (.A(_08541_),
    .B(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__nand2_2 _31095_ (.A(_06051_),
    .B(_06719_),
    .Y(_08544_));
 sky130_fd_sc_hd__o21bai_2 _31096_ (.A1(_08540_),
    .A2(_08543_),
    .B1_N(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__buf_6 _31097_ (.A(_06989_),
    .X(_08546_));
 sky130_fd_sc_hd__nand3b_4 _31098_ (.A_N(_08541_),
    .B(_07333_),
    .C(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand2_1 _31099_ (.A(_08541_),
    .B(_08542_),
    .Y(_08548_));
 sky130_fd_sc_hd__nand3_2 _31100_ (.A(_08547_),
    .B(_08548_),
    .C(_08544_),
    .Y(_08549_));
 sky130_fd_sc_hd__nand2_4 _31101_ (.A(_08545_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__a21o_1 _31102_ (.A1(_08533_),
    .A2(_08539_),
    .B1(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__nand3_4 _31103_ (.A(_08533_),
    .B(_08539_),
    .C(_08550_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_4 _31104_ (.A(_08551_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__o21bai_2 _31105_ (.A1(_08518_),
    .A2(_08521_),
    .B1_N(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__nand3b_4 _31106_ (.A_N(_07982_),
    .B(_08335_),
    .C(_08336_),
    .Y(_08555_));
 sky130_vsdinv _31107_ (.A(_08260_),
    .Y(_08556_));
 sky130_fd_sc_hd__and2_1 _31108_ (.A(_08255_),
    .B(_08263_),
    .X(_08557_));
 sky130_fd_sc_hd__a21oi_4 _31109_ (.A1(_08513_),
    .A2(_08509_),
    .B1(_08516_),
    .Y(_08558_));
 sky130_fd_sc_hd__nor2_1 _31110_ (.A(_08251_),
    .B(_08244_),
    .Y(_08559_));
 sky130_fd_sc_hd__o211a_1 _31111_ (.A1(_08246_),
    .A2(_08559_),
    .B1(_08509_),
    .C1(_08513_),
    .X(_08560_));
 sky130_fd_sc_hd__o22ai_4 _31112_ (.A1(_08556_),
    .A2(_08557_),
    .B1(_08558_),
    .B2(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__o211ai_4 _31113_ (.A1(_08519_),
    .A2(_08520_),
    .B1(_08517_),
    .C1(_08515_),
    .Y(_08562_));
 sky130_fd_sc_hd__nand3_2 _31114_ (.A(_08561_),
    .B(_08562_),
    .C(_08553_),
    .Y(_08563_));
 sky130_fd_sc_hd__nand3_4 _31115_ (.A(_08554_),
    .B(_08555_),
    .C(_08563_),
    .Y(_08564_));
 sky130_vsdinv _31116_ (.A(_08552_),
    .Y(_08565_));
 sky130_vsdinv _31117_ (.A(_08551_),
    .Y(_08566_));
 sky130_fd_sc_hd__o22ai_4 _31118_ (.A1(_08565_),
    .A2(_08566_),
    .B1(_08518_),
    .B2(_08521_),
    .Y(_08567_));
 sky130_fd_sc_hd__nand3b_4 _31119_ (.A_N(_08553_),
    .B(_08561_),
    .C(_08562_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand3_4 _31120_ (.A(_08567_),
    .B(_08339_),
    .C(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__nor2_8 _31121_ (.A(_08300_),
    .B(_08267_),
    .Y(_08570_));
 sky130_fd_sc_hd__nor2_8 _31122_ (.A(_08266_),
    .B(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__nand3_4 _31123_ (.A(_08564_),
    .B(_08569_),
    .C(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__o2bb2ai_4 _31124_ (.A1_N(_08569_),
    .A2_N(_08564_),
    .B1(_08266_),
    .B2(_08570_),
    .Y(_08573_));
 sky130_fd_sc_hd__a21bo_1 _31125_ (.A1(_08323_),
    .A2(_08333_),
    .B1_N(_08324_),
    .X(_08574_));
 sky130_fd_sc_hd__buf_4 _31126_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08575_));
 sky130_fd_sc_hd__and4_4 _31127_ (.A(_19858_),
    .B(_08575_),
    .C(_05313_),
    .D(_05417_),
    .X(_08576_));
 sky130_fd_sc_hd__clkbuf_4 _31128_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08577_));
 sky130_fd_sc_hd__a22o_2 _31129_ (.A1(_19858_),
    .A2(_05417_),
    .B1(_08577_),
    .B2(_05143_),
    .X(_08578_));
 sky130_fd_sc_hd__nand2_2 _31130_ (.A(_19865_),
    .B(_05602_),
    .Y(_08579_));
 sky130_vsdinv _31131_ (.A(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__nand2_1 _31132_ (.A(_08578_),
    .B(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__buf_4 _31133_ (.A(_19857_),
    .X(_08582_));
 sky130_fd_sc_hd__a22oi_4 _31134_ (.A1(_08582_),
    .A2(_05297_),
    .B1(_08577_),
    .B2(_05300_),
    .Y(_08583_));
 sky130_fd_sc_hd__o21ai_2 _31135_ (.A1(_08583_),
    .A2(_08576_),
    .B1(_08579_),
    .Y(_08584_));
 sky130_fd_sc_hd__a31o_1 _31136_ (.A1(_08321_),
    .A2(_19866_),
    .A3(_05181_),
    .B1(_08317_),
    .X(_08585_));
 sky130_fd_sc_hd__o211ai_4 _31137_ (.A1(_08576_),
    .A2(_08581_),
    .B1(_08584_),
    .C1(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__o21ai_2 _31138_ (.A1(_08583_),
    .A2(_08576_),
    .B1(_08580_),
    .Y(_08587_));
 sky130_fd_sc_hd__a21oi_2 _31139_ (.A1(_08319_),
    .A2(_08321_),
    .B1(_08317_),
    .Y(_08588_));
 sky130_fd_sc_hd__buf_4 _31140_ (.A(_19857_),
    .X(_08589_));
 sky130_fd_sc_hd__nand2_1 _31141_ (.A(_08589_),
    .B(_05131_),
    .Y(_08590_));
 sky130_fd_sc_hd__buf_6 _31142_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08591_));
 sky130_fd_sc_hd__buf_6 _31143_ (.A(_08591_),
    .X(_08592_));
 sky130_fd_sc_hd__nand3b_4 _31144_ (.A_N(_08590_),
    .B(_08592_),
    .C(_05179_),
    .Y(_08593_));
 sky130_fd_sc_hd__nand3_2 _31145_ (.A(_08593_),
    .B(_08578_),
    .C(_08579_),
    .Y(_08594_));
 sky130_fd_sc_hd__nand3_4 _31146_ (.A(_08587_),
    .B(_08588_),
    .C(_08594_),
    .Y(_08595_));
 sky130_fd_sc_hd__a22oi_4 _31147_ (.A1(_07482_),
    .A2(_05283_),
    .B1(_07973_),
    .B2(_20162_),
    .Y(_08596_));
 sky130_fd_sc_hd__nand2_2 _31148_ (.A(_07481_),
    .B(_05251_),
    .Y(_08597_));
 sky130_fd_sc_hd__clkbuf_4 _31149_ (.A(\pcpi_mul.rs2[19] ),
    .X(_08598_));
 sky130_fd_sc_hd__nand2_1 _31150_ (.A(_08598_),
    .B(_05392_),
    .Y(_08599_));
 sky130_fd_sc_hd__nor2_1 _31151_ (.A(_08597_),
    .B(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__nand2_2 _31152_ (.A(_07356_),
    .B(_05389_),
    .Y(_08601_));
 sky130_fd_sc_hd__o21bai_2 _31153_ (.A1(_08596_),
    .A2(_08600_),
    .B1_N(_08601_),
    .Y(_08602_));
 sky130_fd_sc_hd__nand3b_4 _31154_ (.A_N(_08597_),
    .B(_08248_),
    .C(_05867_),
    .Y(_08603_));
 sky130_fd_sc_hd__nand2_1 _31155_ (.A(_08597_),
    .B(_08599_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand3_2 _31156_ (.A(_08603_),
    .B(_08604_),
    .C(_08601_),
    .Y(_08605_));
 sky130_fd_sc_hd__nand2_4 _31157_ (.A(_08602_),
    .B(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__a21o_1 _31158_ (.A1(_08586_),
    .A2(_08595_),
    .B1(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__nand3_4 _31159_ (.A(_08586_),
    .B(_08595_),
    .C(_08606_),
    .Y(_08608_));
 sky130_fd_sc_hd__nand3_4 _31160_ (.A(_08574_),
    .B(_08607_),
    .C(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nand2_4 _31161_ (.A(_08607_),
    .B(_08608_),
    .Y(_08610_));
 sky130_fd_sc_hd__a21boi_4 _31162_ (.A1(_08323_),
    .A2(_08333_),
    .B1_N(_08324_),
    .Y(_08611_));
 sky130_fd_sc_hd__nand2_2 _31163_ (.A(_08610_),
    .B(_08611_),
    .Y(_08612_));
 sky130_vsdinv _31164_ (.A(\pcpi_mul.rs2[24] ),
    .Y(_08613_));
 sky130_fd_sc_hd__clkbuf_4 _31165_ (.A(_08613_),
    .X(_08614_));
 sky130_fd_sc_hd__buf_8 _31166_ (.A(net464),
    .X(_08615_));
 sky130_fd_sc_hd__nor2_4 _31167_ (.A(_08615_),
    .B(net449),
    .Y(_08616_));
 sky130_fd_sc_hd__a21oi_4 _31168_ (.A1(_08609_),
    .A2(_08612_),
    .B1(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__and3_2 _31169_ (.A(_08609_),
    .B(_08616_),
    .C(_08612_),
    .X(_08618_));
 sky130_fd_sc_hd__o2bb2ai_4 _31170_ (.A1_N(_08572_),
    .A2_N(_08573_),
    .B1(_08617_),
    .B2(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__nor2_4 _31171_ (.A(_08617_),
    .B(_08618_),
    .Y(_08620_));
 sky130_fd_sc_hd__nand3_4 _31172_ (.A(_08573_),
    .B(_08620_),
    .C(_08572_),
    .Y(_08621_));
 sky130_fd_sc_hd__a21oi_4 _31173_ (.A1(_08619_),
    .A2(_08621_),
    .B1(_08345_),
    .Y(_08622_));
 sky130_fd_sc_hd__and3_2 _31174_ (.A(_08345_),
    .B(_08619_),
    .C(_08621_),
    .X(_08623_));
 sky130_fd_sc_hd__o2bb2ai_4 _31175_ (.A1_N(_08495_),
    .A2_N(_08498_),
    .B1(_08622_),
    .B2(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__and3_4 _31176_ (.A(_08573_),
    .B(_08620_),
    .C(_08572_),
    .X(_08625_));
 sky130_fd_sc_hd__nand2_1 _31177_ (.A(_08345_),
    .B(_08619_),
    .Y(_08626_));
 sky130_fd_sc_hd__nand2_1 _31178_ (.A(_08312_),
    .B(_08341_),
    .Y(_08627_));
 sky130_fd_sc_hd__a21oi_4 _31179_ (.A1(_08573_),
    .A2(_08572_),
    .B1(_08620_),
    .Y(_08628_));
 sky130_fd_sc_hd__o22ai_4 _31180_ (.A1(_08344_),
    .A2(_08627_),
    .B1(_08628_),
    .B2(_08625_),
    .Y(_08629_));
 sky130_fd_sc_hd__o2111ai_4 _31181_ (.A1(_08625_),
    .A2(_08626_),
    .B1(_08629_),
    .C1(_08498_),
    .D1(_08495_),
    .Y(_08630_));
 sky130_fd_sc_hd__nand3_4 _31182_ (.A(_08397_),
    .B(_08624_),
    .C(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand2_1 _31183_ (.A(_08495_),
    .B(_08498_),
    .Y(_08632_));
 sky130_fd_sc_hd__nand3_4 _31184_ (.A(_08345_),
    .B(_08619_),
    .C(_08621_),
    .Y(_08633_));
 sky130_fd_sc_hd__nand3_4 _31185_ (.A(_08632_),
    .B(_08629_),
    .C(_08633_),
    .Y(_08634_));
 sky130_vsdinv _31186_ (.A(_08350_),
    .Y(_08635_));
 sky130_fd_sc_hd__a31oi_4 _31187_ (.A1(_08238_),
    .A2(_08346_),
    .A3(_08240_),
    .B1(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_1 _31188_ (.A(_08629_),
    .B(_08633_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand3_4 _31189_ (.A(_08637_),
    .B(_08495_),
    .C(_08498_),
    .Y(_08638_));
 sky130_fd_sc_hd__nand3_4 _31190_ (.A(_08634_),
    .B(_08636_),
    .C(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__nand2_2 _31191_ (.A(_08239_),
    .B(_08233_),
    .Y(_08640_));
 sky130_fd_sc_hd__nand2_2 _31192_ (.A(_08222_),
    .B(_08217_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand2_2 _31193_ (.A(_08640_),
    .B(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__inv_2 _31194_ (.A(_08642_),
    .Y(_08643_));
 sky130_vsdinv _31195_ (.A(_08641_),
    .Y(_08644_));
 sky130_fd_sc_hd__nand3_4 _31196_ (.A(_08240_),
    .B(_08233_),
    .C(_08644_),
    .Y(_08645_));
 sky130_vsdinv _31197_ (.A(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__o2bb2ai_2 _31198_ (.A1_N(_08631_),
    .A2_N(_08639_),
    .B1(_08643_),
    .B2(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__a21oi_1 _31199_ (.A1(_08358_),
    .A2(_08361_),
    .B1(_08359_),
    .Y(_08648_));
 sky130_fd_sc_hd__o21ai_2 _31200_ (.A1(_08380_),
    .A2(_08648_),
    .B1(_08362_),
    .Y(_08649_));
 sky130_fd_sc_hd__nand2_4 _31201_ (.A(_08642_),
    .B(_08645_),
    .Y(_08650_));
 sky130_vsdinv _31202_ (.A(_08650_),
    .Y(_08651_));
 sky130_fd_sc_hd__nand3_2 _31203_ (.A(_08639_),
    .B(_08651_),
    .C(_08631_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand3_4 _31204_ (.A(_08647_),
    .B(_08649_),
    .C(_08652_),
    .Y(_08653_));
 sky130_vsdinv _31205_ (.A(_08640_),
    .Y(_08654_));
 sky130_fd_sc_hd__nor2_2 _31206_ (.A(_08641_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__nor2_2 _31207_ (.A(_08644_),
    .B(_08640_),
    .Y(_08656_));
 sky130_fd_sc_hd__o2bb2ai_4 _31208_ (.A1_N(_08631_),
    .A2_N(_08639_),
    .B1(_08655_),
    .B2(_08656_),
    .Y(_08657_));
 sky130_fd_sc_hd__a21boi_4 _31209_ (.A1(_08355_),
    .A2(_08366_),
    .B1_N(_08362_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand3_4 _31210_ (.A(_08639_),
    .B(_08631_),
    .C(_08650_),
    .Y(_08659_));
 sky130_fd_sc_hd__nand3_4 _31211_ (.A(_08657_),
    .B(_08658_),
    .C(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__nand2_1 _31212_ (.A(_08653_),
    .B(_08660_),
    .Y(_08661_));
 sky130_vsdinv _31213_ (.A(_08379_),
    .Y(_08662_));
 sky130_fd_sc_hd__nand2_1 _31214_ (.A(_08661_),
    .B(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__a21oi_1 _31215_ (.A1(_08376_),
    .A2(_08381_),
    .B1(_08377_),
    .Y(_08664_));
 sky130_fd_sc_hd__a21oi_2 _31216_ (.A1(_08382_),
    .A2(_08383_),
    .B1(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__nand3_1 _31217_ (.A(_08653_),
    .B(_08660_),
    .C(_08379_),
    .Y(_08666_));
 sky130_fd_sc_hd__nand3_2 _31218_ (.A(_08663_),
    .B(_08665_),
    .C(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__o2bb2ai_1 _31219_ (.A1_N(_08653_),
    .A2_N(_08660_),
    .B1(_08374_),
    .B2(_08372_),
    .Y(_08668_));
 sky130_vsdinv _31220_ (.A(_08368_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand2_1 _31221_ (.A(_08367_),
    .B(_08370_),
    .Y(_08670_));
 sky130_fd_sc_hd__o2bb2ai_2 _31222_ (.A1_N(_08383_),
    .A2_N(_08382_),
    .B1(_08669_),
    .B2(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__nand3_2 _31223_ (.A(_08653_),
    .B(_08660_),
    .C(_08662_),
    .Y(_08672_));
 sky130_fd_sc_hd__nand3_4 _31224_ (.A(_08668_),
    .B(_08671_),
    .C(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__nand2_1 _31225_ (.A(_08667_),
    .B(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__o2111a_2 _31226_ (.A1(_08384_),
    .A2(_08387_),
    .B1(_08132_),
    .C1(_08392_),
    .D1(_08127_),
    .X(_08675_));
 sky130_fd_sc_hd__nand3_4 _31227_ (.A(_08675_),
    .B(_07644_),
    .C(_07884_),
    .Y(_08676_));
 sky130_fd_sc_hd__nor2_8 _31228_ (.A(_07648_),
    .B(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__nor2_1 _31229_ (.A(_08384_),
    .B(_08387_),
    .Y(_08678_));
 sky130_fd_sc_hd__a41o_1 _31230_ (.A1(_08392_),
    .A2(_08130_),
    .A3(_08128_),
    .A4(_08131_),
    .B1(_08678_),
    .X(_08679_));
 sky130_fd_sc_hd__a21oi_4 _31231_ (.A1(_08136_),
    .A2(_08675_),
    .B1(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__o21ai_4 _31232_ (.A1(_08676_),
    .A2(_07651_),
    .B1(_08680_),
    .Y(_08681_));
 sky130_fd_sc_hd__a21oi_4 _31233_ (.A1(_06601_),
    .A2(_08677_),
    .B1(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__nor2_1 _31234_ (.A(_08674_),
    .B(_08682_),
    .Y(_08683_));
 sky130_fd_sc_hd__and2_1 _31235_ (.A(_08682_),
    .B(_08674_),
    .X(_08684_));
 sky130_fd_sc_hd__nor2_2 _31236_ (.A(_08683_),
    .B(_08684_),
    .Y(_02643_));
 sky130_fd_sc_hd__a21oi_2 _31237_ (.A1(_08657_),
    .A2(_08659_),
    .B1(_08658_),
    .Y(_08685_));
 sky130_fd_sc_hd__a21oi_2 _31238_ (.A1(_08662_),
    .A2(_08660_),
    .B1(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand3_1 _31239_ (.A(_08495_),
    .B(_08629_),
    .C(_08497_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_2 _31240_ (.A(_08687_),
    .B(_08633_),
    .Y(_08688_));
 sky130_fd_sc_hd__a22oi_4 _31241_ (.A1(_07294_),
    .A2(_05454_),
    .B1(_07295_),
    .B2(_05827_),
    .Y(_08689_));
 sky130_fd_sc_hd__nand3_4 _31242_ (.A(_07087_),
    .B(_06636_),
    .C(_05453_),
    .Y(_08690_));
 sky130_fd_sc_hd__nor2_8 _31243_ (.A(_06003_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand2_2 _31244_ (.A(_19889_),
    .B(_05825_),
    .Y(_08692_));
 sky130_fd_sc_hd__o21ai_2 _31245_ (.A1(_08689_),
    .A2(_08691_),
    .B1(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__o21ai_4 _31246_ (.A1(_08601_),
    .A2(_08596_),
    .B1(_08603_),
    .Y(_08694_));
 sky130_vsdinv _31247_ (.A(_08692_),
    .Y(_08695_));
 sky130_fd_sc_hd__a22o_2 _31248_ (.A1(_19880_),
    .A2(_06475_),
    .B1(_07755_),
    .B2(_05555_),
    .X(_08696_));
 sky130_fd_sc_hd__o211ai_2 _31249_ (.A1(_06672_),
    .A2(_08690_),
    .B1(_08695_),
    .C1(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__nand3_4 _31250_ (.A(_08693_),
    .B(_08694_),
    .C(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__o21ai_2 _31251_ (.A1(_08689_),
    .A2(_08691_),
    .B1(_08695_),
    .Y(_08699_));
 sky130_fd_sc_hd__o21ai_1 _31252_ (.A1(_08597_),
    .A2(_08599_),
    .B1(_08601_),
    .Y(_08700_));
 sky130_fd_sc_hd__nand2_2 _31253_ (.A(_08700_),
    .B(_08604_),
    .Y(_08701_));
 sky130_fd_sc_hd__o211ai_2 _31254_ (.A1(_06672_),
    .A2(_08690_),
    .B1(_08692_),
    .C1(_08696_),
    .Y(_08702_));
 sky130_fd_sc_hd__nand3_4 _31255_ (.A(_08699_),
    .B(_08701_),
    .C(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__nor2_2 _31256_ (.A(_08505_),
    .B(_08502_),
    .Y(_08704_));
 sky130_fd_sc_hd__o2bb2ai_4 _31257_ (.A1_N(_08698_),
    .A2_N(_08703_),
    .B1(_08500_),
    .B2(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__a21oi_4 _31258_ (.A1(_08506_),
    .A2(_08505_),
    .B1(_08502_),
    .Y(_08706_));
 sky130_fd_sc_hd__nand3b_4 _31259_ (.A_N(_08706_),
    .B(_08698_),
    .C(_08703_),
    .Y(_08707_));
 sky130_fd_sc_hd__nand2_1 _31260_ (.A(_08513_),
    .B(_08516_),
    .Y(_08708_));
 sky130_fd_sc_hd__nand2_4 _31261_ (.A(_08708_),
    .B(_08509_),
    .Y(_08709_));
 sky130_fd_sc_hd__a21oi_4 _31262_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__and3_1 _31263_ (.A(_08504_),
    .B(_08507_),
    .C(_08508_),
    .X(_08711_));
 sky130_fd_sc_hd__nor2_1 _31264_ (.A(_08246_),
    .B(_08559_),
    .Y(_08712_));
 sky130_fd_sc_hd__a31oi_2 _31265_ (.A1(_08510_),
    .A2(_08511_),
    .A3(_08512_),
    .B1(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__o211a_4 _31266_ (.A1(_08711_),
    .A2(_08713_),
    .B1(_08707_),
    .C1(_08705_),
    .X(_08714_));
 sky130_fd_sc_hd__nand2_4 _31267_ (.A(_07785_),
    .B(_06311_),
    .Y(_08715_));
 sky130_fd_sc_hd__a22oi_4 _31268_ (.A1(_07102_),
    .A2(_06695_),
    .B1(_06898_),
    .B2(_06309_),
    .Y(_08716_));
 sky130_fd_sc_hd__nor2_1 _31269_ (.A(_08715_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__nand2_2 _31270_ (.A(_06356_),
    .B(_20141_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand3b_4 _31271_ (.A_N(_08718_),
    .B(_06607_),
    .C(_20138_),
    .Y(_08719_));
 sky130_fd_sc_hd__nand2_2 _31272_ (.A(_08717_),
    .B(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__nand2_2 _31273_ (.A(_08528_),
    .B(_08535_),
    .Y(_08721_));
 sky130_fd_sc_hd__nand2_2 _31274_ (.A(_06545_),
    .B(_07028_),
    .Y(_08722_));
 sky130_fd_sc_hd__nor2_4 _31275_ (.A(_08718_),
    .B(_08722_),
    .Y(_08723_));
 sky130_fd_sc_hd__o21ai_4 _31276_ (.A1(_08716_),
    .A2(_08723_),
    .B1(_08715_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand3_4 _31277_ (.A(_08720_),
    .B(_08721_),
    .C(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__o21bai_2 _31278_ (.A1(_08716_),
    .A2(_08723_),
    .B1_N(_08715_),
    .Y(_08726_));
 sky130_fd_sc_hd__nand2_1 _31279_ (.A(_08718_),
    .B(_08722_),
    .Y(_08727_));
 sky130_fd_sc_hd__nand3_2 _31280_ (.A(_08719_),
    .B(_08727_),
    .C(_08715_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21oi_4 _31281_ (.A1(_08526_),
    .A2(_08527_),
    .B1(_08524_),
    .Y(_08729_));
 sky130_fd_sc_hd__nand3_4 _31282_ (.A(_08726_),
    .B(_08728_),
    .C(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__a22oi_4 _31283_ (.A1(_06627_),
    .A2(_06715_),
    .B1(_06534_),
    .B2(_06813_),
    .Y(_08731_));
 sky130_fd_sc_hd__nand2_1 _31284_ (.A(_06622_),
    .B(_06293_),
    .Y(_08732_));
 sky130_fd_sc_hd__nand2_1 _31285_ (.A(_06044_),
    .B(_06713_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2_2 _31286_ (.A(_08732_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__nand2_2 _31287_ (.A(_06051_),
    .B(_06701_),
    .Y(_08735_));
 sky130_fd_sc_hd__o21bai_2 _31288_ (.A1(_08731_),
    .A2(_08734_),
    .B1_N(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__nand3b_4 _31289_ (.A_N(_08732_),
    .B(_06909_),
    .C(_08151_),
    .Y(_08737_));
 sky130_fd_sc_hd__nand2_1 _31290_ (.A(_08732_),
    .B(_08733_),
    .Y(_08738_));
 sky130_fd_sc_hd__nand3_2 _31291_ (.A(_08737_),
    .B(_08735_),
    .C(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand2_4 _31292_ (.A(_08736_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__a21oi_4 _31293_ (.A1(_08725_),
    .A2(_08730_),
    .B1(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__and3_4 _31294_ (.A(_08725_),
    .B(_08730_),
    .C(_08740_),
    .X(_08742_));
 sky130_fd_sc_hd__nor2_8 _31295_ (.A(_08741_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__o21ai_4 _31296_ (.A1(_08710_),
    .A2(_08714_),
    .B1(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__a21o_1 _31297_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_08709_),
    .X(_08745_));
 sky130_fd_sc_hd__and2_1 _31298_ (.A(_08730_),
    .B(_08740_),
    .X(_08746_));
 sky130_fd_sc_hd__a21o_1 _31299_ (.A1(_08746_),
    .A2(_08725_),
    .B1(_08741_),
    .X(_08747_));
 sky130_fd_sc_hd__nand3_4 _31300_ (.A(_08709_),
    .B(_08705_),
    .C(_08707_),
    .Y(_08748_));
 sky130_fd_sc_hd__nand3_4 _31301_ (.A(_08745_),
    .B(_08747_),
    .C(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand3_4 _31302_ (.A(_08744_),
    .B(_08609_),
    .C(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__o22ai_4 _31303_ (.A1(_08742_),
    .A2(_08741_),
    .B1(_08710_),
    .B2(_08714_),
    .Y(_08751_));
 sky130_fd_sc_hd__nand3_2 _31304_ (.A(_08745_),
    .B(_08743_),
    .C(_08748_),
    .Y(_08752_));
 sky130_fd_sc_hd__nor2_2 _31305_ (.A(_08611_),
    .B(_08610_),
    .Y(_08753_));
 sky130_fd_sc_hd__nand3_4 _31306_ (.A(_08751_),
    .B(_08752_),
    .C(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__o21ai_4 _31307_ (.A1(_08553_),
    .A2(_08518_),
    .B1(_08562_),
    .Y(_08755_));
 sky130_fd_sc_hd__a21oi_4 _31308_ (.A1(_08750_),
    .A2(_08754_),
    .B1(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__and3_1 _31309_ (.A(_08750_),
    .B(_08754_),
    .C(_08755_),
    .X(_08757_));
 sky130_vsdinv _31310_ (.A(_08616_),
    .Y(_08758_));
 sky130_fd_sc_hd__a21oi_4 _31311_ (.A1(_08610_),
    .A2(_08611_),
    .B1(_08758_),
    .Y(_08759_));
 sky130_fd_sc_hd__nand2_1 _31312_ (.A(_08608_),
    .B(_08586_),
    .Y(_08760_));
 sky130_fd_sc_hd__clkbuf_4 _31313_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08761_));
 sky130_fd_sc_hd__and4_4 _31314_ (.A(_08315_),
    .B(_08761_),
    .C(_05456_),
    .D(_05299_),
    .X(_08762_));
 sky130_fd_sc_hd__a22o_1 _31315_ (.A1(_08315_),
    .A2(_05299_),
    .B1(_08761_),
    .B2(_05456_),
    .X(_08763_));
 sky130_fd_sc_hd__nand2_2 _31316_ (.A(\pcpi_mul.rs2[21] ),
    .B(\pcpi_mul.rs1[4] ),
    .Y(_08764_));
 sky130_vsdinv _31317_ (.A(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__nand2_1 _31318_ (.A(_08763_),
    .B(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__o21ai_2 _31319_ (.A1(_08579_),
    .A2(_08583_),
    .B1(_08593_),
    .Y(_08767_));
 sky130_fd_sc_hd__a22oi_4 _31320_ (.A1(_08589_),
    .A2(_05178_),
    .B1(_08575_),
    .B2(_06551_),
    .Y(_08768_));
 sky130_fd_sc_hd__o21ai_2 _31321_ (.A1(_08768_),
    .A2(_08762_),
    .B1(_08764_),
    .Y(_08769_));
 sky130_fd_sc_hd__o211ai_4 _31322_ (.A1(_08762_),
    .A2(_08766_),
    .B1(_08767_),
    .C1(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__o21ai_2 _31323_ (.A1(_08768_),
    .A2(_08762_),
    .B1(_08765_),
    .Y(_08771_));
 sky130_fd_sc_hd__a21oi_4 _31324_ (.A1(_08578_),
    .A2(_08580_),
    .B1(_08576_),
    .Y(_08772_));
 sky130_fd_sc_hd__buf_4 _31325_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08773_));
 sky130_fd_sc_hd__nand2_1 _31326_ (.A(_08773_),
    .B(_20170_),
    .Y(_08774_));
 sky130_fd_sc_hd__clkbuf_4 _31327_ (.A(_08761_),
    .X(_08775_));
 sky130_fd_sc_hd__nand3b_4 _31328_ (.A_N(_08774_),
    .B(_08775_),
    .C(_05245_),
    .Y(_08776_));
 sky130_fd_sc_hd__nand3_2 _31329_ (.A(_08776_),
    .B(_08764_),
    .C(_08763_),
    .Y(_08777_));
 sky130_fd_sc_hd__nand3_4 _31330_ (.A(_08771_),
    .B(_08772_),
    .C(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__buf_4 _31331_ (.A(\pcpi_mul.rs2[20] ),
    .X(_08779_));
 sky130_fd_sc_hd__a22oi_4 _31332_ (.A1(_08779_),
    .A2(_05218_),
    .B1(_07354_),
    .B2(_05389_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand2_2 _31333_ (.A(_07481_),
    .B(_05285_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand2_1 _31334_ (.A(_19872_),
    .B(_05664_),
    .Y(_08782_));
 sky130_fd_sc_hd__nor2_2 _31335_ (.A(_08781_),
    .B(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__nand2_2 _31336_ (.A(_19876_),
    .B(_20155_),
    .Y(_08784_));
 sky130_fd_sc_hd__o21bai_1 _31337_ (.A1(_08780_),
    .A2(_08783_),
    .B1_N(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__nand3b_4 _31338_ (.A_N(_08781_),
    .B(_07973_),
    .C(_05684_),
    .Y(_08786_));
 sky130_fd_sc_hd__nand2_2 _31339_ (.A(_08781_),
    .B(_08782_),
    .Y(_08787_));
 sky130_fd_sc_hd__nand3_1 _31340_ (.A(_08786_),
    .B(_08784_),
    .C(_08787_),
    .Y(_08788_));
 sky130_fd_sc_hd__nand2_2 _31341_ (.A(_08785_),
    .B(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__nand3_2 _31342_ (.A(_08770_),
    .B(_08778_),
    .C(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__nand2_1 _31343_ (.A(_08770_),
    .B(_08778_),
    .Y(_08791_));
 sky130_vsdinv _31344_ (.A(_08789_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand2_1 _31345_ (.A(_08791_),
    .B(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand3_4 _31346_ (.A(_08760_),
    .B(_08790_),
    .C(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__a21boi_2 _31347_ (.A1(_08595_),
    .A2(_08606_),
    .B1_N(_08586_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand2_1 _31348_ (.A(_08791_),
    .B(_08789_),
    .Y(_08796_));
 sky130_fd_sc_hd__nand3_2 _31349_ (.A(_08792_),
    .B(_08778_),
    .C(_08770_),
    .Y(_08797_));
 sky130_fd_sc_hd__nand3_4 _31350_ (.A(_08795_),
    .B(_08796_),
    .C(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__buf_4 _31351_ (.A(\pcpi_mul.rs2[25] ),
    .X(_08799_));
 sky130_fd_sc_hd__clkbuf_4 _31352_ (.A(_08799_),
    .X(_08800_));
 sky130_fd_sc_hd__nand2_4 _31353_ (.A(_08800_),
    .B(_20177_),
    .Y(_08801_));
 sky130_fd_sc_hd__buf_6 _31354_ (.A(\pcpi_mul.rs2[24] ),
    .X(_08802_));
 sky130_fd_sc_hd__nand2_4 _31355_ (.A(_08802_),
    .B(_07901_),
    .Y(_08803_));
 sky130_fd_sc_hd__nor2_8 _31356_ (.A(_08801_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__and2_2 _31357_ (.A(_08801_),
    .B(_08803_),
    .X(_08805_));
 sky130_fd_sc_hd__nor2_8 _31358_ (.A(_08804_),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__a21oi_1 _31359_ (.A1(_08794_),
    .A2(_08798_),
    .B1(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__and3_2 _31360_ (.A(_08794_),
    .B(_08798_),
    .C(_08806_),
    .X(_08808_));
 sky130_fd_sc_hd__o2bb2ai_2 _31361_ (.A1_N(_08609_),
    .A2_N(_08759_),
    .B1(_08807_),
    .B2(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__nand3_4 _31362_ (.A(_08794_),
    .B(_08798_),
    .C(_08806_),
    .Y(_08810_));
 sky130_fd_sc_hd__a21o_1 _31363_ (.A1(_08794_),
    .A2(_08798_),
    .B1(_08806_),
    .X(_08811_));
 sky130_fd_sc_hd__o2111ai_4 _31364_ (.A1(_08610_),
    .A2(_08611_),
    .B1(_08759_),
    .C1(_08810_),
    .D1(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__nand2_2 _31365_ (.A(_08809_),
    .B(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__o21ai_2 _31366_ (.A1(_08756_),
    .A2(_08757_),
    .B1(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__nand3_4 _31367_ (.A(_08750_),
    .B(_08754_),
    .C(_08755_),
    .Y(_08815_));
 sky130_fd_sc_hd__a21o_1 _31368_ (.A1(_08750_),
    .A2(_08754_),
    .B1(_08755_),
    .X(_08816_));
 sky130_fd_sc_hd__nand3b_2 _31369_ (.A_N(_08813_),
    .B(_08815_),
    .C(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__nand3_4 _31370_ (.A(_08625_),
    .B(_08814_),
    .C(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__o21bai_2 _31371_ (.A1(_08756_),
    .A2(_08757_),
    .B1_N(_08813_),
    .Y(_08819_));
 sky130_fd_sc_hd__nand3_2 _31372_ (.A(_08816_),
    .B(_08813_),
    .C(_08815_),
    .Y(_08820_));
 sky130_fd_sc_hd__nand3_4 _31373_ (.A(_08819_),
    .B(_08621_),
    .C(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand2_1 _31374_ (.A(_08818_),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__a22oi_4 _31375_ (.A1(_19911_),
    .A2(_07702_),
    .B1(_05598_),
    .B2(_06993_),
    .Y(_08823_));
 sky130_fd_sc_hd__nand2_4 _31376_ (.A(_07249_),
    .B(_07702_),
    .Y(_08824_));
 sky130_fd_sc_hd__nor2_8 _31377_ (.A(_05860_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__nand2_2 _31378_ (.A(_05865_),
    .B(_20113_),
    .Y(_08826_));
 sky130_fd_sc_hd__o21ai_2 _31379_ (.A1(_08823_),
    .A2(_08825_),
    .B1(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__o21ai_2 _31380_ (.A1(_08544_),
    .A2(_08540_),
    .B1(_08547_),
    .Y(_08828_));
 sky130_vsdinv _31381_ (.A(_08826_),
    .Y(_08829_));
 sky130_fd_sc_hd__a22o_2 _31382_ (.A1(_07660_),
    .A2(_06979_),
    .B1(_05413_),
    .B2(_08042_),
    .X(_08830_));
 sky130_fd_sc_hd__o211ai_4 _31383_ (.A1(_05861_),
    .A2(_08824_),
    .B1(_08829_),
    .C1(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__nand3_4 _31384_ (.A(_08827_),
    .B(_08828_),
    .C(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__o21ai_2 _31385_ (.A1(_08823_),
    .A2(_08825_),
    .B1(_08829_),
    .Y(_08833_));
 sky130_fd_sc_hd__o21ai_1 _31386_ (.A1(_08541_),
    .A2(_08542_),
    .B1(_08544_),
    .Y(_08834_));
 sky130_fd_sc_hd__nand2_2 _31387_ (.A(_08834_),
    .B(_08548_),
    .Y(_08835_));
 sky130_fd_sc_hd__o211ai_4 _31388_ (.A1(_05861_),
    .A2(_08824_),
    .B1(_08826_),
    .C1(_08830_),
    .Y(_08836_));
 sky130_fd_sc_hd__nand3_4 _31389_ (.A(_08833_),
    .B(_08835_),
    .C(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__nor2_4 _31390_ (.A(_08403_),
    .B(_08399_),
    .Y(_08838_));
 sky130_fd_sc_hd__o2bb2ai_4 _31391_ (.A1_N(_08832_),
    .A2_N(_08837_),
    .B1(_08398_),
    .B2(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__nor2_4 _31392_ (.A(_08398_),
    .B(_08838_),
    .Y(_08840_));
 sky130_fd_sc_hd__nand3_4 _31393_ (.A(_08832_),
    .B(_08837_),
    .C(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__nand2_1 _31394_ (.A(_08539_),
    .B(_08550_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_4 _31395_ (.A(_08842_),
    .B(_08533_),
    .Y(_08843_));
 sky130_fd_sc_hd__a21oi_4 _31396_ (.A1(_08839_),
    .A2(_08841_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_vsdinv _31397_ (.A(_08832_),
    .Y(_08845_));
 sky130_fd_sc_hd__nand2_1 _31398_ (.A(_08837_),
    .B(_08840_),
    .Y(_08846_));
 sky130_fd_sc_hd__o211a_1 _31399_ (.A1(_08845_),
    .A2(_08846_),
    .B1(_08839_),
    .C1(_08843_),
    .X(_08847_));
 sky130_fd_sc_hd__nand2_2 _31400_ (.A(_08419_),
    .B(_08406_),
    .Y(_08848_));
 sky130_fd_sc_hd__o21ai_2 _31401_ (.A1(_08844_),
    .A2(_08847_),
    .B1(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__nand2_1 _31402_ (.A(_08425_),
    .B(_08422_),
    .Y(_08850_));
 sky130_fd_sc_hd__nand2_2 _31403_ (.A(_08850_),
    .B(_08424_),
    .Y(_08851_));
 sky130_fd_sc_hd__a21o_1 _31404_ (.A1(_08839_),
    .A2(_08841_),
    .B1(_08843_),
    .X(_08852_));
 sky130_fd_sc_hd__nand3_4 _31405_ (.A(_08843_),
    .B(_08839_),
    .C(_08841_),
    .Y(_08853_));
 sky130_vsdinv _31406_ (.A(_08848_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand3_2 _31407_ (.A(_08852_),
    .B(_08853_),
    .C(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__nand3_4 _31408_ (.A(_08849_),
    .B(_08851_),
    .C(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__o21ai_2 _31409_ (.A1(_08844_),
    .A2(_08847_),
    .B1(_08854_),
    .Y(_08857_));
 sky130_fd_sc_hd__o21ai_2 _31410_ (.A1(_08422_),
    .A2(_08418_),
    .B1(_08425_),
    .Y(_08858_));
 sky130_fd_sc_hd__nand3_2 _31411_ (.A(_08852_),
    .B(_08853_),
    .C(_08848_),
    .Y(_08859_));
 sky130_fd_sc_hd__nand3_4 _31412_ (.A(_08857_),
    .B(_08858_),
    .C(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__a21oi_4 _31413_ (.A1(_08437_),
    .A2(_08439_),
    .B1(_08443_),
    .Y(_08861_));
 sky130_fd_sc_hd__o21ai_2 _31414_ (.A1(_08469_),
    .A2(_08861_),
    .B1(_08444_),
    .Y(_08862_));
 sky130_fd_sc_hd__a21o_1 _31415_ (.A1(_08436_),
    .A2(_08434_),
    .B1(_08432_),
    .X(_08863_));
 sky130_fd_sc_hd__nand2_2 _31416_ (.A(_05311_),
    .B(_07548_),
    .Y(_08864_));
 sky130_fd_sc_hd__nand2_2 _31417_ (.A(_06988_),
    .B(_08196_),
    .Y(_08865_));
 sky130_fd_sc_hd__or2_2 _31418_ (.A(_08864_),
    .B(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__nand2_2 _31419_ (.A(_19937_),
    .B(_20093_),
    .Y(_08867_));
 sky130_vsdinv _31420_ (.A(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__nand2_2 _31421_ (.A(_08864_),
    .B(_08865_),
    .Y(_08869_));
 sky130_fd_sc_hd__nand3_2 _31422_ (.A(_08866_),
    .B(_08868_),
    .C(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__a22oi_4 _31423_ (.A1(_05816_),
    .A2(_07723_),
    .B1(_05978_),
    .B2(_08453_),
    .Y(_08871_));
 sky130_fd_sc_hd__nor2_4 _31424_ (.A(_08864_),
    .B(_08865_),
    .Y(_08872_));
 sky130_fd_sc_hd__o21ai_2 _31425_ (.A1(_08871_),
    .A2(_08872_),
    .B1(_08867_),
    .Y(_08873_));
 sky130_fd_sc_hd__nand3_4 _31426_ (.A(_08863_),
    .B(_08870_),
    .C(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__nand3_2 _31427_ (.A(_08866_),
    .B(_08867_),
    .C(_08869_),
    .Y(_08875_));
 sky130_fd_sc_hd__a21oi_2 _31428_ (.A1(_08436_),
    .A2(_08434_),
    .B1(_08432_),
    .Y(_08876_));
 sky130_fd_sc_hd__o21ai_2 _31429_ (.A1(_08871_),
    .A2(_08872_),
    .B1(_08868_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand3_4 _31430_ (.A(_08875_),
    .B(_08876_),
    .C(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__nand2_1 _31431_ (.A(_08874_),
    .B(_08878_),
    .Y(_08879_));
 sky130_fd_sc_hd__and4_1 _31432_ (.A(_05240_),
    .B(_05242_),
    .C(_20097_),
    .D(_20101_),
    .X(_08880_));
 sky130_fd_sc_hd__clkbuf_4 _31433_ (.A(_08445_),
    .X(_08881_));
 sky130_fd_sc_hd__nand2_1 _31434_ (.A(_05236_),
    .B(_08881_),
    .Y(_08882_));
 sky130_fd_sc_hd__o21a_1 _31435_ (.A1(_05250_),
    .A2(_08435_),
    .B1(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__clkbuf_4 _31436_ (.A(_08447_),
    .X(_08884_));
 sky130_fd_sc_hd__nand2_1 _31437_ (.A(_05692_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__o21ai_1 _31438_ (.A1(_08880_),
    .A2(_08883_),
    .B1(_08885_),
    .Y(_08886_));
 sky130_vsdinv _31439_ (.A(_08885_),
    .Y(_08887_));
 sky130_fd_sc_hd__buf_6 _31440_ (.A(_08435_),
    .X(_08888_));
 sky130_fd_sc_hd__o21ai_2 _31441_ (.A1(_05250_),
    .A2(_08888_),
    .B1(_08882_),
    .Y(_08889_));
 sky130_fd_sc_hd__nand3b_1 _31442_ (.A_N(_08880_),
    .B(_08887_),
    .C(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__nand2_1 _31443_ (.A(_08886_),
    .B(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__nand2_1 _31444_ (.A(_08879_),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__o21ai_1 _31445_ (.A1(_08880_),
    .A2(_08883_),
    .B1(_08887_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand3b_1 _31446_ (.A_N(_08880_),
    .B(_08885_),
    .C(_08889_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand2_2 _31447_ (.A(_08893_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__nand3_2 _31448_ (.A(_08895_),
    .B(_08874_),
    .C(_08878_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand3_4 _31449_ (.A(_08862_),
    .B(_08892_),
    .C(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__nand3_2 _31450_ (.A(_08891_),
    .B(_08874_),
    .C(_08878_),
    .Y(_08898_));
 sky130_fd_sc_hd__nand2_1 _31451_ (.A(_08879_),
    .B(_08895_),
    .Y(_08899_));
 sky130_fd_sc_hd__o2111ai_4 _31452_ (.A1(_08469_),
    .A2(_08861_),
    .B1(_08444_),
    .C1(_08898_),
    .D1(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__nor2_4 _31453_ (.A(_08448_),
    .B(_08451_),
    .Y(_08901_));
 sky130_fd_sc_hd__nor2_8 _31454_ (.A(_08901_),
    .B(_08457_),
    .Y(_08902_));
 sky130_fd_sc_hd__nand3_1 _31455_ (.A(_08897_),
    .B(_08900_),
    .C(_08902_),
    .Y(_08903_));
 sky130_vsdinv _31456_ (.A(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__nand2_2 _31457_ (.A(_08897_),
    .B(_08900_),
    .Y(_08905_));
 sky130_vsdinv _31458_ (.A(_08902_),
    .Y(_08906_));
 sky130_fd_sc_hd__and2_1 _31459_ (.A(_08905_),
    .B(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__o2bb2ai_4 _31460_ (.A1_N(_08856_),
    .A2_N(_08860_),
    .B1(_08904_),
    .B2(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__nand2_1 _31461_ (.A(_08561_),
    .B(_08562_),
    .Y(_08909_));
 sky130_fd_sc_hd__a21oi_2 _31462_ (.A1(_08909_),
    .A2(_08553_),
    .B1(_08555_),
    .Y(_08910_));
 sky130_fd_sc_hd__a22oi_4 _31463_ (.A1(_08910_),
    .A2(_08568_),
    .B1(_08564_),
    .B2(_08571_),
    .Y(_08911_));
 sky130_vsdinv _31464_ (.A(_08897_),
    .Y(_08912_));
 sky130_fd_sc_hd__nand2_1 _31465_ (.A(_08900_),
    .B(_08906_),
    .Y(_08913_));
 sky130_fd_sc_hd__nand2_1 _31466_ (.A(_08905_),
    .B(_08902_),
    .Y(_08914_));
 sky130_fd_sc_hd__o21ai_2 _31467_ (.A1(_08912_),
    .A2(_08913_),
    .B1(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__nand3_4 _31468_ (.A(_08915_),
    .B(_08856_),
    .C(_08860_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand3_4 _31469_ (.A(_08908_),
    .B(_08911_),
    .C(_08916_),
    .Y(_08917_));
 sky130_fd_sc_hd__nor2_1 _31470_ (.A(_08902_),
    .B(_08905_),
    .Y(_08918_));
 sky130_fd_sc_hd__and2_1 _31471_ (.A(_08905_),
    .B(_08902_),
    .X(_08919_));
 sky130_fd_sc_hd__o2bb2ai_1 _31472_ (.A1_N(_08856_),
    .A2_N(_08860_),
    .B1(_08918_),
    .B2(_08919_),
    .Y(_08920_));
 sky130_vsdinv _31473_ (.A(_08568_),
    .Y(_08921_));
 sky130_fd_sc_hd__nand2_1 _31474_ (.A(_08567_),
    .B(_08339_),
    .Y(_08922_));
 sky130_fd_sc_hd__o2bb2ai_2 _31475_ (.A1_N(_08564_),
    .A2_N(_08571_),
    .B1(_08921_),
    .B2(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__nand2_1 _31476_ (.A(_08905_),
    .B(_08906_),
    .Y(_08924_));
 sky130_fd_sc_hd__nand2_1 _31477_ (.A(_08924_),
    .B(_08903_),
    .Y(_08925_));
 sky130_fd_sc_hd__nand3_2 _31478_ (.A(_08925_),
    .B(_08856_),
    .C(_08860_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand3_4 _31479_ (.A(_08920_),
    .B(_08923_),
    .C(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__nor2_2 _31480_ (.A(_08431_),
    .B(_08476_),
    .Y(_08928_));
 sky130_fd_sc_hd__o2bb2ai_4 _31481_ (.A1_N(_08917_),
    .A2_N(_08927_),
    .B1(_08429_),
    .B2(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__o21ai_2 _31482_ (.A1(_08429_),
    .A2(_08483_),
    .B1(_08484_),
    .Y(_08930_));
 sky130_fd_sc_hd__nand3_4 _31483_ (.A(_08927_),
    .B(_08917_),
    .C(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_1 _31484_ (.A(_08929_),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_2 _31485_ (.A(_08822_),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__a21oi_4 _31486_ (.A1(_08908_),
    .A2(_08916_),
    .B1(_08911_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand2_2 _31487_ (.A(_08917_),
    .B(_08930_),
    .Y(_08935_));
 sky130_fd_sc_hd__o2111ai_4 _31488_ (.A1(_08934_),
    .A2(_08935_),
    .B1(_08821_),
    .C1(_08929_),
    .D1(_08818_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand3_4 _31489_ (.A(_08688_),
    .B(_08933_),
    .C(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__a31oi_4 _31490_ (.A1(_08495_),
    .A2(_08629_),
    .A3(_08497_),
    .B1(_08623_),
    .Y(_08938_));
 sky130_fd_sc_hd__nand3_2 _31491_ (.A(_08932_),
    .B(_08821_),
    .C(_08818_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand3_2 _31492_ (.A(_08822_),
    .B(_08929_),
    .C(_08931_),
    .Y(_08940_));
 sky130_fd_sc_hd__nand3_4 _31493_ (.A(_08938_),
    .B(_08939_),
    .C(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand2_1 _31494_ (.A(_08937_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__and2b_2 _31495_ (.A_N(_08473_),
    .B(_08464_),
    .X(_08943_));
 sky130_fd_sc_hd__a21oi_4 _31496_ (.A1(_08497_),
    .A2(_08492_),
    .B1(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__and3_2 _31497_ (.A(_08497_),
    .B(_08492_),
    .C(_08943_),
    .X(_08945_));
 sky130_fd_sc_hd__nor2_8 _31498_ (.A(_08944_),
    .B(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__nand2_1 _31499_ (.A(_08942_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__and2_1 _31500_ (.A(_08633_),
    .B(_08498_),
    .X(_08948_));
 sky130_fd_sc_hd__a21oi_4 _31501_ (.A1(_08493_),
    .A2(_08494_),
    .B1(_08622_),
    .Y(_08949_));
 sky130_fd_sc_hd__a22oi_4 _31502_ (.A1(_08396_),
    .A2(_08350_),
    .B1(_08948_),
    .B2(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__a22oi_4 _31503_ (.A1(_08950_),
    .A2(_08624_),
    .B1(_08639_),
    .B2(_08651_),
    .Y(_08951_));
 sky130_fd_sc_hd__nand3b_2 _31504_ (.A_N(_08946_),
    .B(_08937_),
    .C(_08941_),
    .Y(_08952_));
 sky130_fd_sc_hd__nand3_4 _31505_ (.A(_08947_),
    .B(_08951_),
    .C(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__and3_1 _31506_ (.A(_08397_),
    .B(_08624_),
    .C(_08630_),
    .X(_08954_));
 sky130_fd_sc_hd__a31oi_4 _31507_ (.A1(_08634_),
    .A2(_08636_),
    .A3(_08638_),
    .B1(_08650_),
    .Y(_08955_));
 sky130_fd_sc_hd__nand3_4 _31508_ (.A(_08937_),
    .B(_08941_),
    .C(_08946_),
    .Y(_08956_));
 sky130_fd_sc_hd__o2bb2ai_2 _31509_ (.A1_N(_08941_),
    .A2_N(_08937_),
    .B1(_08944_),
    .B2(_08945_),
    .Y(_08957_));
 sky130_fd_sc_hd__o211ai_4 _31510_ (.A1(_08954_),
    .A2(_08955_),
    .B1(_08956_),
    .C1(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__nand2_1 _31511_ (.A(_08953_),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__nand2_1 _31512_ (.A(_08959_),
    .B(_08642_),
    .Y(_08960_));
 sky130_fd_sc_hd__nand3_4 _31513_ (.A(_08953_),
    .B(_08958_),
    .C(_08643_),
    .Y(_08961_));
 sky130_fd_sc_hd__nand3b_4 _31514_ (.A_N(_08686_),
    .B(_08960_),
    .C(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__nand2_1 _31515_ (.A(_08959_),
    .B(_08643_),
    .Y(_08963_));
 sky130_fd_sc_hd__nand3_1 _31516_ (.A(_08953_),
    .B(_08958_),
    .C(_08642_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand3_2 _31517_ (.A(_08963_),
    .B(_08686_),
    .C(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__and2_2 _31518_ (.A(_08962_),
    .B(_08965_),
    .X(_08966_));
 sky130_fd_sc_hd__o21a_1 _31519_ (.A1(_08674_),
    .A2(_08682_),
    .B1(_08673_),
    .X(_08967_));
 sky130_fd_sc_hd__xnor2_4 _31520_ (.A(_08966_),
    .B(_08967_),
    .Y(_02644_));
 sky130_fd_sc_hd__and2_2 _31521_ (.A(_08913_),
    .B(_08897_),
    .X(_08968_));
 sky130_fd_sc_hd__a21o_2 _31522_ (.A1(_08935_),
    .A2(_08927_),
    .B1(_08968_),
    .X(_08969_));
 sky130_vsdinv _31523_ (.A(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__and2_1 _31524_ (.A(_08935_),
    .B(_08927_),
    .X(_08971_));
 sky130_fd_sc_hd__nand2_2 _31525_ (.A(_08971_),
    .B(_08968_),
    .Y(_08972_));
 sky130_vsdinv _31526_ (.A(_08972_),
    .Y(_08973_));
 sky130_vsdinv _31527_ (.A(_08860_),
    .Y(_08974_));
 sky130_fd_sc_hd__and2_2 _31528_ (.A(_08925_),
    .B(_08856_),
    .X(_08975_));
 sky130_fd_sc_hd__nand2_1 _31529_ (.A(_08750_),
    .B(_08755_),
    .Y(_08976_));
 sky130_fd_sc_hd__nand2_2 _31530_ (.A(_08976_),
    .B(_08754_),
    .Y(_08977_));
 sky130_fd_sc_hd__nand2_1 _31531_ (.A(_08730_),
    .B(_08740_),
    .Y(_08978_));
 sky130_fd_sc_hd__nand2_2 _31532_ (.A(_08978_),
    .B(_08725_),
    .Y(_08979_));
 sky130_fd_sc_hd__a22oi_4 _31533_ (.A1(_19911_),
    .A2(_07249_),
    .B1(_05598_),
    .B2(_08433_),
    .Y(_08980_));
 sky130_fd_sc_hd__and4_2 _31534_ (.A(_06659_),
    .B(_05724_),
    .C(_20113_),
    .D(_07249_),
    .X(_08981_));
 sky130_fd_sc_hd__nand2_2 _31535_ (.A(_05865_),
    .B(_07722_),
    .Y(_08982_));
 sky130_fd_sc_hd__o21ai_2 _31536_ (.A1(_08980_),
    .A2(_08981_),
    .B1(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__nand2_1 _31537_ (.A(_05722_),
    .B(_20117_),
    .Y(_08984_));
 sky130_fd_sc_hd__nand3b_4 _31538_ (.A_N(_08984_),
    .B(_06657_),
    .C(_07564_),
    .Y(_08985_));
 sky130_vsdinv _31539_ (.A(_08982_),
    .Y(_08986_));
 sky130_fd_sc_hd__a22o_1 _31540_ (.A1(_05511_),
    .A2(_06993_),
    .B1(_05598_),
    .B2(_08433_),
    .X(_08987_));
 sky130_fd_sc_hd__nand3_2 _31541_ (.A(_08985_),
    .B(_08986_),
    .C(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__o21ai_2 _31542_ (.A1(_08735_),
    .A2(_08731_),
    .B1(_08737_),
    .Y(_08989_));
 sky130_fd_sc_hd__nand3_4 _31543_ (.A(_08983_),
    .B(_08988_),
    .C(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__o21ai_2 _31544_ (.A1(_08980_),
    .A2(_08981_),
    .B1(_08986_),
    .Y(_08991_));
 sky130_fd_sc_hd__nand3_2 _31545_ (.A(_08985_),
    .B(_08982_),
    .C(_08987_),
    .Y(_08992_));
 sky130_vsdinv _31546_ (.A(_08735_),
    .Y(_08993_));
 sky130_fd_sc_hd__a21oi_2 _31547_ (.A1(_08993_),
    .A2(_08738_),
    .B1(_08734_),
    .Y(_08994_));
 sky130_fd_sc_hd__nand3_4 _31548_ (.A(_08991_),
    .B(_08992_),
    .C(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__nor2_4 _31549_ (.A(_08829_),
    .B(_08825_),
    .Y(_08996_));
 sky130_fd_sc_hd__o2bb2ai_4 _31550_ (.A1_N(_08990_),
    .A2_N(_08995_),
    .B1(_08823_),
    .B2(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__nor2_4 _31551_ (.A(_08823_),
    .B(_08996_),
    .Y(_08998_));
 sky130_fd_sc_hd__nand3_4 _31552_ (.A(_08990_),
    .B(_08995_),
    .C(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__nand3_4 _31553_ (.A(_08979_),
    .B(_08997_),
    .C(_08999_),
    .Y(_09000_));
 sky130_vsdinv _31554_ (.A(_08730_),
    .Y(_09001_));
 sky130_fd_sc_hd__a31oi_4 _31555_ (.A1(_08721_),
    .A2(_08720_),
    .A3(_08724_),
    .B1(_08740_),
    .Y(_09002_));
 sky130_fd_sc_hd__a21oi_4 _31556_ (.A1(_08990_),
    .A2(_08995_),
    .B1(_08998_),
    .Y(_09003_));
 sky130_fd_sc_hd__nor2_1 _31557_ (.A(_08826_),
    .B(_08823_),
    .Y(_09004_));
 sky130_fd_sc_hd__o211a_1 _31558_ (.A1(_08825_),
    .A2(_09004_),
    .B1(_08990_),
    .C1(_08995_),
    .X(_09005_));
 sky130_fd_sc_hd__o22ai_4 _31559_ (.A1(_09001_),
    .A2(_09002_),
    .B1(_09003_),
    .B2(_09005_),
    .Y(_09006_));
 sky130_vsdinv _31560_ (.A(_08837_),
    .Y(_09007_));
 sky130_fd_sc_hd__nor2_1 _31561_ (.A(_08840_),
    .B(_08845_),
    .Y(_09008_));
 sky130_fd_sc_hd__o2bb2ai_1 _31562_ (.A1_N(_09000_),
    .A2_N(_09006_),
    .B1(_09007_),
    .B2(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__and2_1 _31563_ (.A(_08837_),
    .B(_08840_),
    .X(_09010_));
 sky130_fd_sc_hd__nor2_4 _31564_ (.A(_08845_),
    .B(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand3b_2 _31565_ (.A_N(_09011_),
    .B(_09006_),
    .C(_09000_),
    .Y(_09012_));
 sky130_fd_sc_hd__o21ai_2 _31566_ (.A1(_08854_),
    .A2(_08844_),
    .B1(_08853_),
    .Y(_09013_));
 sky130_fd_sc_hd__nand3_4 _31567_ (.A(_09009_),
    .B(_09012_),
    .C(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__o2bb2ai_1 _31568_ (.A1_N(_09000_),
    .A2_N(_09006_),
    .B1(_08845_),
    .B2(_09010_),
    .Y(_09015_));
 sky130_fd_sc_hd__nand2_1 _31569_ (.A(_08853_),
    .B(_08854_),
    .Y(_09016_));
 sky130_fd_sc_hd__nand2_2 _31570_ (.A(_09016_),
    .B(_08852_),
    .Y(_09017_));
 sky130_fd_sc_hd__nand3_2 _31571_ (.A(_09006_),
    .B(_09000_),
    .C(_09011_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand3_4 _31572_ (.A(_09015_),
    .B(_09017_),
    .C(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__nand2_2 _31573_ (.A(_05376_),
    .B(_08196_),
    .Y(_09020_));
 sky130_fd_sc_hd__nand2_2 _31574_ (.A(_05211_),
    .B(_08036_),
    .Y(_09021_));
 sky130_fd_sc_hd__or2_4 _31575_ (.A(_09020_),
    .B(_09021_),
    .X(_09022_));
 sky130_fd_sc_hd__a22oi_4 _31576_ (.A1(_06986_),
    .A2(_08196_),
    .B1(_06988_),
    .B2(_08447_),
    .Y(_09023_));
 sky130_vsdinv _31577_ (.A(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__clkbuf_4 _31578_ (.A(\pcpi_mul.rs1[26] ),
    .X(_09025_));
 sky130_fd_sc_hd__nand2_4 _31579_ (.A(_05192_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__nand3_2 _31580_ (.A(_09022_),
    .B(_09024_),
    .C(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__a21oi_2 _31581_ (.A1(_08868_),
    .A2(_08869_),
    .B1(_08872_),
    .Y(_09028_));
 sky130_fd_sc_hd__nor2_2 _31582_ (.A(_09020_),
    .B(_09021_),
    .Y(_09029_));
 sky130_vsdinv _31583_ (.A(_09026_),
    .Y(_09030_));
 sky130_fd_sc_hd__o21ai_2 _31584_ (.A1(_09023_),
    .A2(_09029_),
    .B1(_09030_),
    .Y(_09031_));
 sky130_fd_sc_hd__nand3_4 _31585_ (.A(_09027_),
    .B(_09028_),
    .C(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__nand3_2 _31586_ (.A(_09022_),
    .B(_09024_),
    .C(_09030_),
    .Y(_09033_));
 sky130_fd_sc_hd__a21o_1 _31587_ (.A1(_08868_),
    .A2(_08869_),
    .B1(_08872_),
    .X(_09034_));
 sky130_fd_sc_hd__o21ai_2 _31588_ (.A1(_09023_),
    .A2(_09029_),
    .B1(_09026_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand3_4 _31589_ (.A(_09033_),
    .B(_09034_),
    .C(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__clkbuf_4 _31590_ (.A(\pcpi_mul.rs1[25] ),
    .X(_09037_));
 sky130_fd_sc_hd__buf_4 _31591_ (.A(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__nand2_1 _31592_ (.A(_05139_),
    .B(_20097_),
    .Y(_09039_));
 sky130_fd_sc_hd__a21o_1 _31593_ (.A1(_19934_),
    .A2(_09038_),
    .B1(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__buf_4 _31594_ (.A(_20096_),
    .X(_09041_));
 sky130_fd_sc_hd__nand2_1 _31595_ (.A(_05141_),
    .B(_20093_),
    .Y(_09042_));
 sky130_fd_sc_hd__a21o_1 _31596_ (.A1(_06314_),
    .A2(_09041_),
    .B1(_09042_),
    .X(_09043_));
 sky130_fd_sc_hd__buf_6 _31597_ (.A(_20101_),
    .X(_09044_));
 sky130_fd_sc_hd__nand2_2 _31598_ (.A(_19928_),
    .B(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__a21oi_4 _31599_ (.A1(_09040_),
    .A2(_09043_),
    .B1(_09045_),
    .Y(_09046_));
 sky130_vsdinv _31600_ (.A(_08445_),
    .Y(_09047_));
 sky130_fd_sc_hd__o211a_2 _31601_ (.A1(_05186_),
    .A2(_09047_),
    .B1(_09043_),
    .C1(_09040_),
    .X(_09048_));
 sky130_fd_sc_hd__nor2_8 _31602_ (.A(_09046_),
    .B(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__a21o_1 _31603_ (.A1(_09032_),
    .A2(_09036_),
    .B1(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__nand3_4 _31604_ (.A(_09049_),
    .B(_09036_),
    .C(_09032_),
    .Y(_09051_));
 sky130_fd_sc_hd__nand2_1 _31605_ (.A(_08895_),
    .B(_08878_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand2_2 _31606_ (.A(_09052_),
    .B(_08874_),
    .Y(_09053_));
 sky130_fd_sc_hd__a21o_2 _31607_ (.A1(_09050_),
    .A2(_09051_),
    .B1(_09053_),
    .X(_09054_));
 sky130_fd_sc_hd__nand3_4 _31608_ (.A(_09050_),
    .B(_09053_),
    .C(_09051_),
    .Y(_09055_));
 sky130_fd_sc_hd__a21o_2 _31609_ (.A1(_08889_),
    .A2(_08887_),
    .B1(_08880_),
    .X(_09056_));
 sky130_fd_sc_hd__a21oi_4 _31610_ (.A1(_09054_),
    .A2(_09055_),
    .B1(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__and3_1 _31611_ (.A(_09054_),
    .B(_09056_),
    .C(_09055_),
    .X(_09058_));
 sky130_fd_sc_hd__o2bb2ai_4 _31612_ (.A1_N(_09014_),
    .A2_N(_09019_),
    .B1(_09057_),
    .B2(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__a21oi_1 _31613_ (.A1(_09050_),
    .A2(_09051_),
    .B1(_09053_),
    .Y(_09060_));
 sky130_vsdinv _31614_ (.A(_09036_),
    .Y(_09061_));
 sky130_fd_sc_hd__nand2_1 _31615_ (.A(_09049_),
    .B(_09032_),
    .Y(_09062_));
 sky130_fd_sc_hd__o211a_1 _31616_ (.A1(_09061_),
    .A2(_09062_),
    .B1(_09053_),
    .C1(_09050_),
    .X(_09063_));
 sky130_fd_sc_hd__o21ai_2 _31617_ (.A1(_09060_),
    .A2(_09063_),
    .B1(_09056_),
    .Y(_09064_));
 sky130_fd_sc_hd__nand3b_2 _31618_ (.A_N(_09056_),
    .B(_09054_),
    .C(_09055_),
    .Y(_09065_));
 sky130_fd_sc_hd__nand2_4 _31619_ (.A(_09064_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__nand3_4 _31620_ (.A(_09066_),
    .B(_09014_),
    .C(_09019_),
    .Y(_09067_));
 sky130_fd_sc_hd__nand3_4 _31621_ (.A(_08977_),
    .B(_09059_),
    .C(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__nand2_2 _31622_ (.A(_09059_),
    .B(_09067_),
    .Y(_09069_));
 sky130_fd_sc_hd__o21a_1 _31623_ (.A1(_08553_),
    .A2(_08518_),
    .B1(_08562_),
    .X(_09070_));
 sky130_fd_sc_hd__a31oi_4 _31624_ (.A1(_08744_),
    .A2(_08749_),
    .A3(_08609_),
    .B1(_09070_),
    .Y(_09071_));
 sky130_vsdinv _31625_ (.A(_08754_),
    .Y(_09072_));
 sky130_fd_sc_hd__nor2_2 _31626_ (.A(_09071_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__nand2_1 _31627_ (.A(_09069_),
    .B(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__o211ai_4 _31628_ (.A1(_08974_),
    .A2(_08975_),
    .B1(_09068_),
    .C1(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__a21oi_2 _31629_ (.A1(_09059_),
    .A2(_09067_),
    .B1(_08977_),
    .Y(_09076_));
 sky130_fd_sc_hd__o211a_2 _31630_ (.A1(_09072_),
    .A2(_09071_),
    .B1(_09067_),
    .C1(_09059_),
    .X(_09077_));
 sky130_fd_sc_hd__nor2_2 _31631_ (.A(_08974_),
    .B(_08975_),
    .Y(_09078_));
 sky130_fd_sc_hd__o21ai_4 _31632_ (.A1(_09076_),
    .A2(_09077_),
    .B1(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__nand2_4 _31633_ (.A(_08698_),
    .B(_08706_),
    .Y(_09080_));
 sky130_fd_sc_hd__a22oi_4 _31634_ (.A1(_06927_),
    .A2(_05689_),
    .B1(_06925_),
    .B2(_20145_),
    .Y(_09081_));
 sky130_fd_sc_hd__nand3_4 _31635_ (.A(_07753_),
    .B(_19885_),
    .C(_05554_),
    .Y(_09082_));
 sky130_fd_sc_hd__nor2_4 _31636_ (.A(_06287_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__nand2_2 _31637_ (.A(_19889_),
    .B(_06152_),
    .Y(_09084_));
 sky130_vsdinv _31638_ (.A(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__o21ai_2 _31639_ (.A1(_09081_),
    .A2(_09083_),
    .B1(_09085_),
    .Y(_09086_));
 sky130_vsdinv _31640_ (.A(_08784_),
    .Y(_09087_));
 sky130_fd_sc_hd__a21oi_4 _31641_ (.A1(_09087_),
    .A2(_08787_),
    .B1(_08783_),
    .Y(_09088_));
 sky130_fd_sc_hd__a22o_2 _31642_ (.A1(_19880_),
    .A2(_05689_),
    .B1(_07755_),
    .B2(_05822_),
    .X(_09089_));
 sky130_fd_sc_hd__o211ai_4 _31643_ (.A1(_06287_),
    .A2(_09082_),
    .B1(_09084_),
    .C1(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__nand3_4 _31644_ (.A(_09086_),
    .B(_09088_),
    .C(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__o21ai_2 _31645_ (.A1(_09081_),
    .A2(_09083_),
    .B1(_09084_),
    .Y(_09092_));
 sky130_fd_sc_hd__o21ai_4 _31646_ (.A1(_08784_),
    .A2(_08780_),
    .B1(_08786_),
    .Y(_09093_));
 sky130_fd_sc_hd__o211ai_4 _31647_ (.A1(_06297_),
    .A2(_09082_),
    .B1(_09085_),
    .C1(_09089_),
    .Y(_09094_));
 sky130_fd_sc_hd__nand3_4 _31648_ (.A(_09092_),
    .B(_09093_),
    .C(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__nor2_2 _31649_ (.A(_08695_),
    .B(_08691_),
    .Y(_09096_));
 sky130_fd_sc_hd__o2bb2ai_4 _31650_ (.A1_N(_09091_),
    .A2_N(_09095_),
    .B1(_08689_),
    .B2(_09096_),
    .Y(_09097_));
 sky130_fd_sc_hd__a21oi_4 _31651_ (.A1(_08696_),
    .A2(_08695_),
    .B1(_08691_),
    .Y(_09098_));
 sky130_vsdinv _31652_ (.A(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__nand3_4 _31653_ (.A(_09091_),
    .B(_09095_),
    .C(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__a22oi_4 _31654_ (.A1(_08703_),
    .A2(_09080_),
    .B1(_09097_),
    .B2(_09100_),
    .Y(_09101_));
 sky130_fd_sc_hd__a21oi_4 _31655_ (.A1(_09091_),
    .A2(_09095_),
    .B1(_09099_),
    .Y(_09102_));
 sky130_fd_sc_hd__nand3_4 _31656_ (.A(_09100_),
    .B(_08703_),
    .C(_09080_),
    .Y(_09103_));
 sky130_fd_sc_hd__nor2_8 _31657_ (.A(_09102_),
    .B(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__a22oi_4 _31658_ (.A1(_07922_),
    .A2(_06696_),
    .B1(_06207_),
    .B2(_07661_),
    .Y(_09105_));
 sky130_fd_sc_hd__and4_2 _31659_ (.A(_07102_),
    .B(_19895_),
    .C(_06142_),
    .D(_07028_),
    .X(_09106_));
 sky130_fd_sc_hd__nand2_2 _31660_ (.A(\pcpi_mul.rs2[12] ),
    .B(_20132_),
    .Y(_09107_));
 sky130_fd_sc_hd__o21ai_2 _31661_ (.A1(_09105_),
    .A2(_09106_),
    .B1(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__nand2_1 _31662_ (.A(_06543_),
    .B(_05985_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand3b_4 _31663_ (.A_N(_09109_),
    .B(_06895_),
    .C(_07503_),
    .Y(_09110_));
 sky130_vsdinv _31664_ (.A(_09107_),
    .Y(_09111_));
 sky130_fd_sc_hd__a22o_2 _31665_ (.A1(_07922_),
    .A2(_06309_),
    .B1(_06898_),
    .B2(_06311_),
    .X(_09112_));
 sky130_fd_sc_hd__nand3_2 _31666_ (.A(_09110_),
    .B(_09111_),
    .C(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__o21ai_2 _31667_ (.A1(_08715_),
    .A2(_08716_),
    .B1(_08719_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand3_4 _31668_ (.A(_09108_),
    .B(_09113_),
    .C(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__o21ai_2 _31669_ (.A1(_09105_),
    .A2(_09106_),
    .B1(_09111_),
    .Y(_09116_));
 sky130_fd_sc_hd__nand3_2 _31670_ (.A(_09110_),
    .B(_09107_),
    .C(_09112_),
    .Y(_09117_));
 sky130_fd_sc_hd__o21ai_1 _31671_ (.A1(_08718_),
    .A2(_08722_),
    .B1(_08715_),
    .Y(_09118_));
 sky130_fd_sc_hd__nand2_1 _31672_ (.A(_09118_),
    .B(_08727_),
    .Y(_09119_));
 sky130_fd_sc_hd__nand3_4 _31673_ (.A(_09116_),
    .B(_09117_),
    .C(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__a22oi_4 _31674_ (.A1(_06627_),
    .A2(_06813_),
    .B1(_06631_),
    .B2(_06816_),
    .Y(_09121_));
 sky130_fd_sc_hd__nand2_2 _31675_ (.A(_06622_),
    .B(_20128_),
    .Y(_09122_));
 sky130_fd_sc_hd__nand2_2 _31676_ (.A(_06044_),
    .B(_06701_),
    .Y(_09123_));
 sky130_fd_sc_hd__nor2_4 _31677_ (.A(_09122_),
    .B(_09123_),
    .Y(_09124_));
 sky130_fd_sc_hd__nand2_2 _31678_ (.A(_05952_),
    .B(_07251_),
    .Y(_09125_));
 sky130_fd_sc_hd__o21bai_2 _31679_ (.A1(_09121_),
    .A2(_09124_),
    .B1_N(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand3b_4 _31680_ (.A_N(_09122_),
    .B(_05657_),
    .C(_07709_),
    .Y(_09127_));
 sky130_fd_sc_hd__nand2_2 _31681_ (.A(_09122_),
    .B(_09123_),
    .Y(_09128_));
 sky130_fd_sc_hd__nand3_2 _31682_ (.A(_09127_),
    .B(_09125_),
    .C(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__nand2_4 _31683_ (.A(_09126_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__a21oi_4 _31684_ (.A1(_09115_),
    .A2(_09120_),
    .B1(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__and3_2 _31685_ (.A(_09120_),
    .B(_09115_),
    .C(_09130_),
    .X(_09132_));
 sky130_fd_sc_hd__nor2_8 _31686_ (.A(_09131_),
    .B(_09132_),
    .Y(_09133_));
 sky130_fd_sc_hd__o21ai_2 _31687_ (.A1(_09101_),
    .A2(_09104_),
    .B1(_09133_),
    .Y(_09134_));
 sky130_fd_sc_hd__a22o_2 _31688_ (.A1(_08703_),
    .A2(_09080_),
    .B1(_09097_),
    .B2(_09100_),
    .X(_09135_));
 sky130_fd_sc_hd__and2_1 _31689_ (.A(_09120_),
    .B(_09130_),
    .X(_09136_));
 sky130_fd_sc_hd__a21o_1 _31690_ (.A1(_09136_),
    .A2(_09115_),
    .B1(_09131_),
    .X(_09137_));
 sky130_fd_sc_hd__and3_1 _31691_ (.A(_09092_),
    .B(_09093_),
    .C(_09094_),
    .X(_09138_));
 sky130_fd_sc_hd__nand2_2 _31692_ (.A(_09091_),
    .B(_09099_),
    .Y(_09139_));
 sky130_fd_sc_hd__o2111ai_4 _31693_ (.A1(_09138_),
    .A2(_09139_),
    .B1(_08703_),
    .C1(_09097_),
    .D1(_09080_),
    .Y(_09140_));
 sky130_fd_sc_hd__nand3_2 _31694_ (.A(_09135_),
    .B(_09137_),
    .C(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__nand3_4 _31695_ (.A(_09134_),
    .B(_08794_),
    .C(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__o22ai_4 _31696_ (.A1(_09132_),
    .A2(_09131_),
    .B1(_09101_),
    .B2(_09104_),
    .Y(_09143_));
 sky130_fd_sc_hd__nand3_2 _31697_ (.A(_09135_),
    .B(_09140_),
    .C(_09133_),
    .Y(_09144_));
 sky130_vsdinv _31698_ (.A(_08794_),
    .Y(_09145_));
 sky130_fd_sc_hd__nand3_4 _31699_ (.A(_09143_),
    .B(_09144_),
    .C(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__nor2_8 _31700_ (.A(_08743_),
    .B(_08714_),
    .Y(_09147_));
 sky130_fd_sc_hd__nor2_8 _31701_ (.A(_08710_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__nand3_4 _31702_ (.A(_09142_),
    .B(_09146_),
    .C(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__o2bb2ai_4 _31703_ (.A1_N(_09146_),
    .A2_N(_09142_),
    .B1(_08710_),
    .B2(_09147_),
    .Y(_09150_));
 sky130_fd_sc_hd__a22oi_4 _31704_ (.A1(_08315_),
    .A2(_05456_),
    .B1(_08761_),
    .B2(_20164_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_2 _31705_ (.A(\pcpi_mul.rs2[23] ),
    .B(\pcpi_mul.rs1[3] ),
    .Y(_09152_));
 sky130_fd_sc_hd__nand2_2 _31706_ (.A(_08761_),
    .B(_05243_),
    .Y(_09153_));
 sky130_fd_sc_hd__nor2_4 _31707_ (.A(_09152_),
    .B(_09153_),
    .Y(_09154_));
 sky130_fd_sc_hd__nand2_2 _31708_ (.A(\pcpi_mul.rs2[21] ),
    .B(_20161_),
    .Y(_09155_));
 sky130_fd_sc_hd__o21ai_2 _31709_ (.A1(_09151_),
    .A2(_09154_),
    .B1(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__nand3b_4 _31710_ (.A_N(_09152_),
    .B(_08591_),
    .C(_05460_),
    .Y(_09157_));
 sky130_vsdinv _31711_ (.A(_09155_),
    .Y(_09158_));
 sky130_fd_sc_hd__nand2_2 _31712_ (.A(_09152_),
    .B(_09153_),
    .Y(_09159_));
 sky130_fd_sc_hd__nand3_2 _31713_ (.A(_09157_),
    .B(_09158_),
    .C(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__o21ai_2 _31714_ (.A1(_08764_),
    .A2(_08768_),
    .B1(_08776_),
    .Y(_09161_));
 sky130_fd_sc_hd__nand3_4 _31715_ (.A(_09156_),
    .B(_09160_),
    .C(_09161_),
    .Y(_09162_));
 sky130_fd_sc_hd__a21oi_2 _31716_ (.A1(_08763_),
    .A2(_08765_),
    .B1(_08762_),
    .Y(_09163_));
 sky130_fd_sc_hd__o21ai_2 _31717_ (.A1(_09151_),
    .A2(_09154_),
    .B1(_09158_),
    .Y(_09164_));
 sky130_fd_sc_hd__nand3_2 _31718_ (.A(_09157_),
    .B(_09155_),
    .C(_09159_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand3_4 _31719_ (.A(_09163_),
    .B(_09164_),
    .C(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__a22oi_4 _31720_ (.A1(_07481_),
    .A2(_05294_),
    .B1(_19872_),
    .B2(_05372_),
    .Y(_09167_));
 sky130_fd_sc_hd__nand2_2 _31721_ (.A(\pcpi_mul.rs2[20] ),
    .B(\pcpi_mul.rs1[6] ),
    .Y(_09168_));
 sky130_fd_sc_hd__nand2_1 _31722_ (.A(\pcpi_mul.rs2[19] ),
    .B(_05372_),
    .Y(_09169_));
 sky130_fd_sc_hd__nor2_2 _31723_ (.A(_09168_),
    .B(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__nand2_2 _31724_ (.A(\pcpi_mul.rs2[18] ),
    .B(\pcpi_mul.rs1[8] ),
    .Y(_09171_));
 sky130_fd_sc_hd__o21a_1 _31725_ (.A1(_09167_),
    .A2(_09170_),
    .B1(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__nand3b_4 _31726_ (.A_N(_09168_),
    .B(_07827_),
    .C(_20155_),
    .Y(_09173_));
 sky130_vsdinv _31727_ (.A(_09171_),
    .Y(_09174_));
 sky130_fd_sc_hd__nand2_1 _31728_ (.A(_09168_),
    .B(_09169_),
    .Y(_09175_));
 sky130_fd_sc_hd__and3_1 _31729_ (.A(_09173_),
    .B(_09174_),
    .C(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__o2bb2ai_4 _31730_ (.A1_N(_09162_),
    .A2_N(_09166_),
    .B1(_09172_),
    .B2(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__o21ai_1 _31731_ (.A1(_09167_),
    .A2(_09170_),
    .B1(_09174_),
    .Y(_09178_));
 sky130_fd_sc_hd__nand3_1 _31732_ (.A(_09173_),
    .B(_09171_),
    .C(_09175_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_2 _31733_ (.A(_09178_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__nand3_4 _31734_ (.A(_09166_),
    .B(_09162_),
    .C(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__nand2_1 _31735_ (.A(_08778_),
    .B(_08789_),
    .Y(_09182_));
 sky130_fd_sc_hd__nand2_4 _31736_ (.A(_09182_),
    .B(_08770_),
    .Y(_09183_));
 sky130_fd_sc_hd__a21oi_2 _31737_ (.A1(_09177_),
    .A2(_09181_),
    .B1(_09183_),
    .Y(_09184_));
 sky130_vsdinv _31738_ (.A(_09162_),
    .Y(_09185_));
 sky130_fd_sc_hd__nand2_2 _31739_ (.A(_09166_),
    .B(_09180_),
    .Y(_09186_));
 sky130_fd_sc_hd__o211a_1 _31740_ (.A1(_09185_),
    .A2(_09186_),
    .B1(_09177_),
    .C1(_09183_),
    .X(_09187_));
 sky130_vsdinv _31741_ (.A(_08804_),
    .Y(_09188_));
 sky130_fd_sc_hd__nand2_4 _31742_ (.A(_08799_),
    .B(_05145_),
    .Y(_09189_));
 sky130_fd_sc_hd__nand2_4 _31743_ (.A(_19846_),
    .B(_20176_),
    .Y(_09190_));
 sky130_fd_sc_hd__nor2_4 _31744_ (.A(_09189_),
    .B(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__and2_1 _31745_ (.A(_09189_),
    .B(_09190_),
    .X(_09192_));
 sky130_fd_sc_hd__nor2_8 _31746_ (.A(_08613_),
    .B(_05126_),
    .Y(_09193_));
 sky130_fd_sc_hd__o21bai_2 _31747_ (.A1(_09191_),
    .A2(_09192_),
    .B1_N(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_2 _31748_ (.A(_09189_),
    .B(_09190_),
    .Y(_09195_));
 sky130_fd_sc_hd__nand3b_2 _31749_ (.A_N(_09191_),
    .B(_09195_),
    .C(_09193_),
    .Y(_09196_));
 sky130_fd_sc_hd__nand2_4 _31750_ (.A(_09194_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__nor2_8 _31751_ (.A(_09188_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand2_1 _31752_ (.A(_09197_),
    .B(_09188_),
    .Y(_09199_));
 sky130_fd_sc_hd__or2b_4 _31753_ (.A(_09198_),
    .B_N(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__o21ai_4 _31754_ (.A1(_09184_),
    .A2(_09187_),
    .B1(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__a21o_1 _31755_ (.A1(_09177_),
    .A2(_09181_),
    .B1(_09183_),
    .X(_09202_));
 sky130_fd_sc_hd__nand3_4 _31756_ (.A(_09183_),
    .B(_09177_),
    .C(_09181_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand3b_4 _31757_ (.A_N(_09200_),
    .B(_09202_),
    .C(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__a21oi_2 _31758_ (.A1(_09201_),
    .A2(_09204_),
    .B1(_08808_),
    .Y(_09205_));
 sky130_fd_sc_hd__nand3_4 _31759_ (.A(_08808_),
    .B(_09201_),
    .C(_09204_),
    .Y(_09206_));
 sky130_vsdinv _31760_ (.A(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__o2bb2ai_4 _31761_ (.A1_N(_09149_),
    .A2_N(_09150_),
    .B1(_09205_),
    .B2(_09207_),
    .Y(_09208_));
 sky130_vsdinv _31762_ (.A(_09204_),
    .Y(_09209_));
 sky130_fd_sc_hd__nand2_1 _31763_ (.A(_08808_),
    .B(_09201_),
    .Y(_09210_));
 sky130_fd_sc_hd__nand2_2 _31764_ (.A(_09201_),
    .B(_09204_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_4 _31765_ (.A(_09211_),
    .B(_08810_),
    .Y(_09212_));
 sky130_fd_sc_hd__o2111ai_4 _31766_ (.A1(_09209_),
    .A2(_09210_),
    .B1(_09212_),
    .C1(_09149_),
    .D1(_09150_),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_2 _31767_ (.A(_08815_),
    .B(_08809_),
    .Y(_09214_));
 sky130_fd_sc_hd__o21ai_4 _31768_ (.A1(_08756_),
    .A2(_09214_),
    .B1(_08812_),
    .Y(_09215_));
 sky130_fd_sc_hd__a21oi_2 _31769_ (.A1(_09208_),
    .A2(_09213_),
    .B1(_09215_),
    .Y(_09216_));
 sky130_fd_sc_hd__a21oi_4 _31770_ (.A1(_09142_),
    .A2(_09146_),
    .B1(_09148_),
    .Y(_09217_));
 sky130_fd_sc_hd__nand3_4 _31771_ (.A(_09149_),
    .B(_09212_),
    .C(_09206_),
    .Y(_09218_));
 sky130_fd_sc_hd__o211a_2 _31772_ (.A1(_09217_),
    .A2(_09218_),
    .B1(_09208_),
    .C1(_09215_),
    .X(_09219_));
 sky130_fd_sc_hd__o2bb2ai_4 _31773_ (.A1_N(_09075_),
    .A2_N(_09079_),
    .B1(_09216_),
    .B2(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__o2bb2ai_4 _31774_ (.A1_N(_09073_),
    .A2_N(_09069_),
    .B1(_08974_),
    .B2(_08975_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand3_4 _31775_ (.A(_09215_),
    .B(_09208_),
    .C(_09213_),
    .Y(_09222_));
 sky130_fd_sc_hd__a22oi_4 _31776_ (.A1(_09212_),
    .A2(_09206_),
    .B1(_09150_),
    .B2(_09149_),
    .Y(_09223_));
 sky130_fd_sc_hd__nor2_2 _31777_ (.A(_09217_),
    .B(_09218_),
    .Y(_09224_));
 sky130_fd_sc_hd__o21a_1 _31778_ (.A1(_08756_),
    .A2(_09214_),
    .B1(_08812_),
    .X(_09225_));
 sky130_fd_sc_hd__o21ai_4 _31779_ (.A1(_09223_),
    .A2(_09224_),
    .B1(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__o2111ai_4 _31780_ (.A1(_09077_),
    .A2(_09221_),
    .B1(_09222_),
    .C1(_09226_),
    .D1(_09079_),
    .Y(_09227_));
 sky130_fd_sc_hd__nand3_1 _31781_ (.A(_08929_),
    .B(_08821_),
    .C(_08931_),
    .Y(_09228_));
 sky130_fd_sc_hd__nand2_2 _31782_ (.A(_09228_),
    .B(_08818_),
    .Y(_09229_));
 sky130_fd_sc_hd__a21oi_4 _31783_ (.A1(_09220_),
    .A2(_09227_),
    .B1(_09229_),
    .Y(_09230_));
 sky130_vsdinv _31784_ (.A(_08818_),
    .Y(_09231_));
 sky130_fd_sc_hd__o211a_1 _31785_ (.A1(_08934_),
    .A2(_08935_),
    .B1(_08821_),
    .C1(_08929_),
    .X(_09232_));
 sky130_fd_sc_hd__o211a_2 _31786_ (.A1(_09231_),
    .A2(_09232_),
    .B1(_09220_),
    .C1(_09227_),
    .X(_09233_));
 sky130_fd_sc_hd__o22ai_4 _31787_ (.A1(_08970_),
    .A2(_08973_),
    .B1(_09230_),
    .B2(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_4 _31788_ (.A(_08972_),
    .B(_08969_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand2_1 _31789_ (.A(_09220_),
    .B(_09227_),
    .Y(_09236_));
 sky130_fd_sc_hd__nor2_1 _31790_ (.A(_09231_),
    .B(_09232_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_2 _31791_ (.A(_09236_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__nand3_4 _31792_ (.A(_09220_),
    .B(_09227_),
    .C(_09229_),
    .Y(_09239_));
 sky130_fd_sc_hd__nand3b_4 _31793_ (.A_N(_09235_),
    .B(_09238_),
    .C(_09239_),
    .Y(_09240_));
 sky130_vsdinv _31794_ (.A(_08933_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand2_1 _31795_ (.A(_08688_),
    .B(_08936_),
    .Y(_09242_));
 sky130_fd_sc_hd__o2bb2ai_2 _31796_ (.A1_N(_08941_),
    .A2_N(_08946_),
    .B1(_09241_),
    .B2(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__nand3_4 _31797_ (.A(_09234_),
    .B(_09240_),
    .C(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__o21bai_2 _31798_ (.A1(_09230_),
    .A2(_09233_),
    .B1_N(_09235_),
    .Y(_09245_));
 sky130_fd_sc_hd__a21boi_4 _31799_ (.A1(_08941_),
    .A2(_08946_),
    .B1_N(_08937_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand3_4 _31800_ (.A(_09238_),
    .B(_09239_),
    .C(_09235_),
    .Y(_09247_));
 sky130_fd_sc_hd__nand3_4 _31801_ (.A(_09245_),
    .B(_09246_),
    .C(_09247_),
    .Y(_09248_));
 sky130_fd_sc_hd__and2_1 _31802_ (.A(_08498_),
    .B(_08492_),
    .X(_09249_));
 sky130_fd_sc_hd__o2bb2ai_2 _31803_ (.A1_N(_09244_),
    .A2_N(_09248_),
    .B1(_08943_),
    .B2(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand3_2 _31804_ (.A(_09248_),
    .B(_09244_),
    .C(_08944_),
    .Y(_09251_));
 sky130_fd_sc_hd__o21ai_1 _31805_ (.A1(_08954_),
    .A2(_08955_),
    .B1(_08957_),
    .Y(_09252_));
 sky130_vsdinv _31806_ (.A(_08956_),
    .Y(_09253_));
 sky130_fd_sc_hd__o2bb2ai_2 _31807_ (.A1_N(_08643_),
    .A2_N(_08953_),
    .B1(_09252_),
    .B2(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__a21oi_4 _31808_ (.A1(_09250_),
    .A2(_09251_),
    .B1(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__and3_1 _31809_ (.A(_09245_),
    .B(_09246_),
    .C(_09247_),
    .X(_09256_));
 sky130_fd_sc_hd__nand2_1 _31810_ (.A(_09244_),
    .B(_08944_),
    .Y(_09257_));
 sky130_fd_sc_hd__o211a_2 _31811_ (.A1(_09256_),
    .A2(_09257_),
    .B1(_09254_),
    .C1(_09250_),
    .X(_09258_));
 sky130_fd_sc_hd__nor2_8 _31812_ (.A(_09255_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__a21boi_4 _31813_ (.A1(_08962_),
    .A2(_08673_),
    .B1_N(_08965_),
    .Y(_09260_));
 sky130_fd_sc_hd__a21oi_1 _31814_ (.A1(_08953_),
    .A2(_08958_),
    .B1(_08643_),
    .Y(_09261_));
 sky130_fd_sc_hd__a31oi_1 _31815_ (.A1(_08657_),
    .A2(_08658_),
    .A3(_08659_),
    .B1(_08379_),
    .Y(_09262_));
 sky130_fd_sc_hd__o21ai_1 _31816_ (.A1(_08685_),
    .A2(_09262_),
    .B1(_08961_),
    .Y(_09263_));
 sky130_fd_sc_hd__o2111a_2 _31817_ (.A1(_09261_),
    .A2(_09263_),
    .B1(_08673_),
    .C1(_08667_),
    .D1(_08965_),
    .X(_09264_));
 sky130_fd_sc_hd__and2b_2 _31818_ (.A_N(_08682_),
    .B(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__nor2_8 _31819_ (.A(_09260_),
    .B(_09265_),
    .Y(_09266_));
 sky130_fd_sc_hd__xnor2_4 _31820_ (.A(_09259_),
    .B(_09266_),
    .Y(_02645_));
 sky130_fd_sc_hd__a31oi_4 _31821_ (.A1(_09079_),
    .A2(_09226_),
    .A3(_09075_),
    .B1(_09219_),
    .Y(_09267_));
 sky130_fd_sc_hd__a22oi_4 _31822_ (.A1(_08773_),
    .A2(_20164_),
    .B1(_08591_),
    .B2(_05289_),
    .Y(_09268_));
 sky130_vsdinv _31823_ (.A(_20161_),
    .Y(_09269_));
 sky130_fd_sc_hd__nand3_4 _31824_ (.A(_19857_),
    .B(\pcpi_mul.rs2[22] ),
    .C(_05243_),
    .Y(_09270_));
 sky130_fd_sc_hd__nor2_4 _31825_ (.A(_09269_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__nand2_4 _31826_ (.A(\pcpi_mul.rs2[21] ),
    .B(_05294_),
    .Y(_09272_));
 sky130_fd_sc_hd__o21ai_2 _31827_ (.A1(_09268_),
    .A2(_09271_),
    .B1(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__o21ai_2 _31828_ (.A1(_09155_),
    .A2(_09151_),
    .B1(_09157_),
    .Y(_09274_));
 sky130_fd_sc_hd__buf_6 _31829_ (.A(_09269_),
    .X(_09275_));
 sky130_vsdinv _31830_ (.A(_09272_),
    .Y(_09276_));
 sky130_fd_sc_hd__a22o_2 _31831_ (.A1(_08315_),
    .A2(_20164_),
    .B1(_19862_),
    .B2(_05480_),
    .X(_09277_));
 sky130_fd_sc_hd__o211ai_4 _31832_ (.A1(_09275_),
    .A2(_09270_),
    .B1(_09276_),
    .C1(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__nand3_4 _31833_ (.A(_09273_),
    .B(_09274_),
    .C(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__o21ai_2 _31834_ (.A1(_09268_),
    .A2(_09271_),
    .B1(_09276_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21oi_2 _31835_ (.A1(_09158_),
    .A2(_09159_),
    .B1(_09154_),
    .Y(_09281_));
 sky130_fd_sc_hd__o211ai_4 _31836_ (.A1(_09275_),
    .A2(_09270_),
    .B1(_09272_),
    .C1(_09277_),
    .Y(_09282_));
 sky130_fd_sc_hd__nand3_4 _31837_ (.A(_09280_),
    .B(_09281_),
    .C(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__a22oi_4 _31838_ (.A1(_08779_),
    .A2(_05472_),
    .B1(_08598_),
    .B2(_05571_),
    .Y(_09284_));
 sky130_fd_sc_hd__nand3_4 _31839_ (.A(_07481_),
    .B(\pcpi_mul.rs2[19] ),
    .C(_05372_),
    .Y(_09285_));
 sky130_fd_sc_hd__nor2_4 _31840_ (.A(_08242_),
    .B(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__nand2_4 _31841_ (.A(\pcpi_mul.rs2[18] ),
    .B(_20148_),
    .Y(_09287_));
 sky130_fd_sc_hd__o21a_1 _31842_ (.A1(_09284_),
    .A2(_09286_),
    .B1(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__nor3_4 _31843_ (.A(_09287_),
    .B(_09284_),
    .C(_09286_),
    .Y(_09289_));
 sky130_fd_sc_hd__o2bb2ai_4 _31844_ (.A1_N(_09279_),
    .A2_N(_09283_),
    .B1(_09288_),
    .B2(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__a22o_1 _31845_ (.A1(_08779_),
    .A2(_05696_),
    .B1(_08598_),
    .B2(_05571_),
    .X(_09291_));
 sky130_fd_sc_hd__nand3b_1 _31846_ (.A_N(_09286_),
    .B(_09291_),
    .C(_09287_),
    .Y(_09292_));
 sky130_vsdinv _31847_ (.A(_09287_),
    .Y(_09293_));
 sky130_fd_sc_hd__o21ai_1 _31848_ (.A1(_09284_),
    .A2(_09286_),
    .B1(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__nand2_1 _31849_ (.A(_09292_),
    .B(_09294_),
    .Y(_09295_));
 sky130_fd_sc_hd__nand3_4 _31850_ (.A(_09295_),
    .B(_09283_),
    .C(_09279_),
    .Y(_09296_));
 sky130_fd_sc_hd__a21oi_4 _31851_ (.A1(_09290_),
    .A2(_09296_),
    .B1(_09198_),
    .Y(_09297_));
 sky130_fd_sc_hd__nand3_4 _31852_ (.A(_09290_),
    .B(_09198_),
    .C(_09296_),
    .Y(_09298_));
 sky130_fd_sc_hd__nand2_4 _31853_ (.A(_09186_),
    .B(_09162_),
    .Y(_09299_));
 sky130_fd_sc_hd__nand2_1 _31854_ (.A(_09298_),
    .B(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__nor2_4 _31855_ (.A(_09297_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__o2bb2ai_4 _31856_ (.A1_N(_09296_),
    .A2_N(_09290_),
    .B1(_09188_),
    .B2(_09197_),
    .Y(_09302_));
 sky130_fd_sc_hd__a21oi_4 _31857_ (.A1(_09302_),
    .A2(_09298_),
    .B1(_09299_),
    .Y(_09303_));
 sky130_fd_sc_hd__a21oi_4 _31858_ (.A1(_09193_),
    .A2(_09195_),
    .B1(_09191_),
    .Y(_09304_));
 sky130_fd_sc_hd__nand2_4 _31859_ (.A(_19846_),
    .B(\pcpi_mul.rs1[1] ),
    .Y(_09305_));
 sky130_fd_sc_hd__nand2_4 _31860_ (.A(_08799_),
    .B(_05125_),
    .Y(_09306_));
 sky130_fd_sc_hd__nor2_8 _31861_ (.A(_09305_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__nand2_4 _31862_ (.A(_09305_),
    .B(_09306_),
    .Y(_09308_));
 sky130_vsdinv _31863_ (.A(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__nor2_8 _31864_ (.A(_08613_),
    .B(_05369_),
    .Y(_09310_));
 sky130_vsdinv _31865_ (.A(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__o21ai_2 _31866_ (.A1(_09307_),
    .A2(_09309_),
    .B1(_09311_),
    .Y(_09312_));
 sky130_vsdinv _31867_ (.A(_09307_),
    .Y(_09313_));
 sky130_fd_sc_hd__nand3_4 _31868_ (.A(_09313_),
    .B(_09310_),
    .C(_09308_),
    .Y(_09314_));
 sky130_fd_sc_hd__nand3b_4 _31869_ (.A_N(_09304_),
    .B(_09312_),
    .C(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__nand3_2 _31870_ (.A(_09311_),
    .B(_09313_),
    .C(_09308_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ai_2 _31871_ (.A1(_09307_),
    .A2(_09309_),
    .B1(_09310_),
    .Y(_09317_));
 sky130_fd_sc_hd__nand3_4 _31872_ (.A(_09316_),
    .B(_09317_),
    .C(_09304_),
    .Y(_09318_));
 sky130_fd_sc_hd__nand2_1 _31873_ (.A(_09315_),
    .B(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__buf_8 _31874_ (.A(\pcpi_mul.rs2[27] ),
    .X(_09320_));
 sky130_fd_sc_hd__inv_4 _31875_ (.A(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__nor2_2 _31876_ (.A(_09321_),
    .B(net449),
    .Y(_09322_));
 sky130_vsdinv _31877_ (.A(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__nand2_1 _31878_ (.A(_09319_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nand3_4 _31879_ (.A(_09315_),
    .B(_09318_),
    .C(_09322_),
    .Y(_09325_));
 sky130_fd_sc_hd__nand2_2 _31880_ (.A(_09324_),
    .B(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__o21ai_4 _31881_ (.A1(_09301_),
    .A2(_09303_),
    .B1(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__and3_1 _31882_ (.A(_09290_),
    .B(_09198_),
    .C(_09296_),
    .X(_09328_));
 sky130_vsdinv _31883_ (.A(_09299_),
    .Y(_09329_));
 sky130_fd_sc_hd__o21ai_2 _31884_ (.A1(_09297_),
    .A2(_09328_),
    .B1(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__nand3_4 _31885_ (.A(_09302_),
    .B(_09298_),
    .C(_09299_),
    .Y(_09331_));
 sky130_vsdinv _31886_ (.A(_09326_),
    .Y(_09332_));
 sky130_fd_sc_hd__nand3_4 _31887_ (.A(_09330_),
    .B(_09331_),
    .C(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__a21oi_4 _31888_ (.A1(_09327_),
    .A2(_09333_),
    .B1(_09209_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _31889_ (.A(_09330_),
    .B(_09332_),
    .Y(_09335_));
 sky130_fd_sc_hd__o211a_2 _31890_ (.A1(_09301_),
    .A2(_09335_),
    .B1(_09209_),
    .C1(_09327_),
    .X(_09336_));
 sky130_fd_sc_hd__nand2_2 _31891_ (.A(_06356_),
    .B(_06441_),
    .Y(_09337_));
 sky130_fd_sc_hd__nand2_2 _31892_ (.A(\pcpi_mul.rs2[13] ),
    .B(_06293_),
    .Y(_09338_));
 sky130_fd_sc_hd__or2_1 _31893_ (.A(_09337_),
    .B(_09338_),
    .X(_09339_));
 sky130_fd_sc_hd__nand2_2 _31894_ (.A(\pcpi_mul.rs2[12] ),
    .B(_20128_),
    .Y(_09340_));
 sky130_vsdinv _31895_ (.A(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__nand2_2 _31896_ (.A(_09337_),
    .B(_09338_),
    .Y(_09342_));
 sky130_fd_sc_hd__nand3_2 _31897_ (.A(_09339_),
    .B(_09341_),
    .C(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__o21ai_2 _31898_ (.A1(_09107_),
    .A2(_09105_),
    .B1(_09110_),
    .Y(_09344_));
 sky130_fd_sc_hd__a22oi_4 _31899_ (.A1(_07922_),
    .A2(_06438_),
    .B1(_06607_),
    .B2(_06437_),
    .Y(_09345_));
 sky130_fd_sc_hd__nor2_4 _31900_ (.A(_09337_),
    .B(_09338_),
    .Y(_09346_));
 sky130_fd_sc_hd__o21ai_2 _31901_ (.A1(_09345_),
    .A2(_09346_),
    .B1(_09340_),
    .Y(_09347_));
 sky130_fd_sc_hd__nand3_2 _31902_ (.A(_09343_),
    .B(_09344_),
    .C(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__nand3_2 _31903_ (.A(_09339_),
    .B(_09340_),
    .C(_09342_),
    .Y(_09349_));
 sky130_fd_sc_hd__a21oi_4 _31904_ (.A1(_09112_),
    .A2(_09111_),
    .B1(_09106_),
    .Y(_09350_));
 sky130_fd_sc_hd__o21ai_2 _31905_ (.A1(_09345_),
    .A2(_09346_),
    .B1(_09341_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand3_4 _31906_ (.A(_09349_),
    .B(_09350_),
    .C(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_2 _31907_ (.A(_06117_),
    .B(_20125_),
    .Y(_09353_));
 sky130_fd_sc_hd__nand2_2 _31908_ (.A(_05656_),
    .B(_20122_),
    .Y(_09354_));
 sky130_fd_sc_hd__or2_1 _31909_ (.A(_09353_),
    .B(_09354_),
    .X(_09355_));
 sky130_fd_sc_hd__nand2_1 _31910_ (.A(_06051_),
    .B(_06993_),
    .Y(_09356_));
 sky130_fd_sc_hd__nand2_2 _31911_ (.A(_09353_),
    .B(_09354_),
    .Y(_09357_));
 sky130_fd_sc_hd__nand3_2 _31912_ (.A(_09355_),
    .B(_09356_),
    .C(_09357_),
    .Y(_09358_));
 sky130_fd_sc_hd__a22oi_2 _31913_ (.A1(_06630_),
    .A2(_08142_),
    .B1(_06909_),
    .B2(_07567_),
    .Y(_09359_));
 sky130_fd_sc_hd__nor2_4 _31914_ (.A(_09353_),
    .B(_09354_),
    .Y(_09360_));
 sky130_vsdinv _31915_ (.A(_09356_),
    .Y(_09361_));
 sky130_fd_sc_hd__o21ai_2 _31916_ (.A1(_09359_),
    .A2(_09360_),
    .B1(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__nand2_4 _31917_ (.A(_09358_),
    .B(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__nand3_1 _31918_ (.A(_09348_),
    .B(_09352_),
    .C(_09363_),
    .Y(_09364_));
 sky130_vsdinv _31919_ (.A(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__nand2_1 _31920_ (.A(_09348_),
    .B(_09352_),
    .Y(_09366_));
 sky130_vsdinv _31921_ (.A(_09363_),
    .Y(_09367_));
 sky130_fd_sc_hd__and2_1 _31922_ (.A(_09366_),
    .B(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__a22oi_4 _31923_ (.A1(_07753_),
    .A2(_05825_),
    .B1(_06636_),
    .B2(_06152_),
    .Y(_09369_));
 sky130_fd_sc_hd__and4_4 _31924_ (.A(\pcpi_mul.rs2[17] ),
    .B(_19885_),
    .C(_06152_),
    .D(_20144_),
    .X(_09370_));
 sky130_fd_sc_hd__o22ai_4 _31925_ (.A1(_06528_),
    .A2(_06445_),
    .B1(_09369_),
    .B2(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__o21ai_2 _31926_ (.A1(_09171_),
    .A2(_09167_),
    .B1(_09173_),
    .Y(_09372_));
 sky130_fd_sc_hd__nand2_2 _31927_ (.A(\pcpi_mul.rs2[15] ),
    .B(\pcpi_mul.rs1[12] ),
    .Y(_09373_));
 sky130_fd_sc_hd__a41oi_2 _31928_ (.A1(_06927_),
    .A2(_07089_),
    .A3(_05998_),
    .A4(_05670_),
    .B1(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__a22o_1 _31929_ (.A1(_07087_),
    .A2(_05825_),
    .B1(_07089_),
    .B2(_20141_),
    .X(_09375_));
 sky130_fd_sc_hd__nand2_2 _31930_ (.A(_09374_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand3_4 _31931_ (.A(_09371_),
    .B(_09372_),
    .C(_09376_),
    .Y(_09377_));
 sky130_vsdinv _31932_ (.A(_09373_),
    .Y(_09378_));
 sky130_fd_sc_hd__o21ai_2 _31933_ (.A1(_09369_),
    .A2(_09370_),
    .B1(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__nand2_1 _31934_ (.A(_07753_),
    .B(_05825_),
    .Y(_09380_));
 sky130_fd_sc_hd__nand3b_2 _31935_ (.A_N(_09380_),
    .B(_07755_),
    .C(_06695_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand3_4 _31936_ (.A(_09381_),
    .B(_09373_),
    .C(_09375_),
    .Y(_09382_));
 sky130_fd_sc_hd__a21oi_2 _31937_ (.A1(_09174_),
    .A2(_09175_),
    .B1(_09170_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand3_4 _31938_ (.A(_09379_),
    .B(_09382_),
    .C(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__nor2_4 _31939_ (.A(_09085_),
    .B(_09083_),
    .Y(_09385_));
 sky130_fd_sc_hd__o2bb2ai_4 _31940_ (.A1_N(_09377_),
    .A2_N(_09384_),
    .B1(_09081_),
    .B2(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__nor2_2 _31941_ (.A(_09081_),
    .B(_09385_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand3_4 _31942_ (.A(_09384_),
    .B(_09377_),
    .C(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__nand2_4 _31943_ (.A(_09139_),
    .B(_09095_),
    .Y(_09389_));
 sky130_fd_sc_hd__a21oi_4 _31944_ (.A1(_09386_),
    .A2(_09388_),
    .B1(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__a31oi_2 _31945_ (.A1(_09086_),
    .A2(_09088_),
    .A3(_09090_),
    .B1(_09098_),
    .Y(_09391_));
 sky130_fd_sc_hd__o211a_4 _31946_ (.A1(_09138_),
    .A2(_09391_),
    .B1(_09388_),
    .C1(_09386_),
    .X(_09392_));
 sky130_fd_sc_hd__o22ai_2 _31947_ (.A1(_09365_),
    .A2(_09368_),
    .B1(_09390_),
    .B2(_09392_),
    .Y(_09393_));
 sky130_fd_sc_hd__a21o_2 _31948_ (.A1(_09386_),
    .A2(_09388_),
    .B1(_09389_),
    .X(_09394_));
 sky130_fd_sc_hd__nand3_2 _31949_ (.A(_09367_),
    .B(_09352_),
    .C(_09348_),
    .Y(_09395_));
 sky130_fd_sc_hd__nand2_1 _31950_ (.A(_09366_),
    .B(_09363_),
    .Y(_09396_));
 sky130_fd_sc_hd__nand2_4 _31951_ (.A(_09395_),
    .B(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__nand3_4 _31952_ (.A(_09389_),
    .B(_09386_),
    .C(_09388_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand3_1 _31953_ (.A(_09394_),
    .B(_09397_),
    .C(_09398_),
    .Y(_09399_));
 sky130_fd_sc_hd__nand3_2 _31954_ (.A(_09393_),
    .B(_09187_),
    .C(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__buf_2 _31955_ (.A(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__o21ai_4 _31956_ (.A1(_09390_),
    .A2(_09392_),
    .B1(_09397_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand2_1 _31957_ (.A(_09366_),
    .B(_09367_),
    .Y(_09403_));
 sky130_fd_sc_hd__nand2_1 _31958_ (.A(_09403_),
    .B(_09364_),
    .Y(_09404_));
 sky130_fd_sc_hd__nand3_4 _31959_ (.A(_09394_),
    .B(_09404_),
    .C(_09398_),
    .Y(_09405_));
 sky130_fd_sc_hd__a21oi_4 _31960_ (.A1(_09135_),
    .A2(_09133_),
    .B1(_09104_),
    .Y(_09406_));
 sky130_fd_sc_hd__a31oi_4 _31961_ (.A1(_09402_),
    .A2(_09405_),
    .A3(_09203_),
    .B1(_09406_),
    .Y(_09407_));
 sky130_fd_sc_hd__nand3_4 _31962_ (.A(_09402_),
    .B(_09203_),
    .C(_09405_),
    .Y(_09408_));
 sky130_vsdinv _31963_ (.A(_09406_),
    .Y(_09409_));
 sky130_fd_sc_hd__a21oi_4 _31964_ (.A1(_09408_),
    .A2(_09401_),
    .B1(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__a21oi_1 _31965_ (.A1(_09401_),
    .A2(_09407_),
    .B1(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__o21ai_2 _31966_ (.A1(_09334_),
    .A2(_09336_),
    .B1(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__a31oi_4 _31967_ (.A1(_09150_),
    .A2(_09212_),
    .A3(_09149_),
    .B1(_09207_),
    .Y(_09413_));
 sky130_fd_sc_hd__nor2_1 _31968_ (.A(_09133_),
    .B(_09104_),
    .Y(_09414_));
 sky130_fd_sc_hd__o2bb2ai_2 _31969_ (.A1_N(_09400_),
    .A2_N(_09408_),
    .B1(_09101_),
    .B2(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__nand3_1 _31970_ (.A(_09409_),
    .B(_09401_),
    .C(_09408_),
    .Y(_09416_));
 sky130_fd_sc_hd__nand2_2 _31971_ (.A(_09415_),
    .B(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__nand2_1 _31972_ (.A(_09202_),
    .B(_09203_),
    .Y(_09418_));
 sky130_fd_sc_hd__o2bb2ai_2 _31973_ (.A1_N(_09333_),
    .A2_N(_09327_),
    .B1(_09418_),
    .B2(_09200_),
    .Y(_09419_));
 sky130_fd_sc_hd__nand3_4 _31974_ (.A(_09327_),
    .B(_09209_),
    .C(_09333_),
    .Y(_09420_));
 sky130_fd_sc_hd__nand3_2 _31975_ (.A(_09417_),
    .B(_09419_),
    .C(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand3_4 _31976_ (.A(_09412_),
    .B(_09413_),
    .C(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__nor2_1 _31977_ (.A(_09101_),
    .B(_09137_),
    .Y(_09423_));
 sky130_fd_sc_hd__o211a_1 _31978_ (.A1(_09104_),
    .A2(_09423_),
    .B1(_09401_),
    .C1(_09408_),
    .X(_09424_));
 sky130_fd_sc_hd__o22ai_4 _31979_ (.A1(_09424_),
    .A2(_09410_),
    .B1(_09334_),
    .B2(_09336_),
    .Y(_09425_));
 sky130_vsdinv _31980_ (.A(_09401_),
    .Y(_09426_));
 sky130_fd_sc_hd__nand2_2 _31981_ (.A(_09409_),
    .B(_09408_),
    .Y(_09427_));
 sky130_fd_sc_hd__o2111ai_4 _31982_ (.A1(_09426_),
    .A2(_09427_),
    .B1(_09420_),
    .C1(_09415_),
    .D1(_09419_),
    .Y(_09428_));
 sky130_fd_sc_hd__o22ai_4 _31983_ (.A1(_08810_),
    .A2(_09211_),
    .B1(_09217_),
    .B2(_09218_),
    .Y(_09429_));
 sky130_fd_sc_hd__nand3_4 _31984_ (.A(_09425_),
    .B(_09428_),
    .C(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__nand2_1 _31985_ (.A(_09422_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__a22oi_4 _31986_ (.A1(_06659_),
    .A2(_20113_),
    .B1(_05598_),
    .B2(_07722_),
    .Y(_09432_));
 sky130_vsdinv _31987_ (.A(\pcpi_mul.rs1[20] ),
    .Y(_09433_));
 sky130_fd_sc_hd__nand3_4 _31988_ (.A(_05501_),
    .B(_19914_),
    .C(_07232_),
    .Y(_09434_));
 sky130_fd_sc_hd__nor2_4 _31989_ (.A(_09433_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__nand2_2 _31990_ (.A(_05865_),
    .B(\pcpi_mul.rs1[21] ),
    .Y(_09436_));
 sky130_fd_sc_hd__o21ai_2 _31991_ (.A1(_09432_),
    .A2(_09435_),
    .B1(_09436_),
    .Y(_09437_));
 sky130_vsdinv _31992_ (.A(_09436_),
    .Y(_09438_));
 sky130_fd_sc_hd__a22o_2 _31993_ (.A1(_05511_),
    .A2(_08433_),
    .B1(_06840_),
    .B2(_07722_),
    .X(_09439_));
 sky130_fd_sc_hd__o211ai_4 _31994_ (.A1(_09433_),
    .A2(_09434_),
    .B1(_09438_),
    .C1(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__o21ai_4 _31995_ (.A1(_09125_),
    .A2(_09121_),
    .B1(_09127_),
    .Y(_09441_));
 sky130_fd_sc_hd__nand3_4 _31996_ (.A(_09437_),
    .B(_09440_),
    .C(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__clkbuf_8 _31997_ (.A(_06979_),
    .X(_09443_));
 sky130_fd_sc_hd__a31oi_4 _31998_ (.A1(_09128_),
    .A2(_06052_),
    .A3(_09443_),
    .B1(_09124_),
    .Y(_09444_));
 sky130_fd_sc_hd__o21ai_2 _31999_ (.A1(_09432_),
    .A2(_09435_),
    .B1(_09438_),
    .Y(_09445_));
 sky130_fd_sc_hd__o211ai_4 _32000_ (.A1(_09433_),
    .A2(_09434_),
    .B1(_09436_),
    .C1(_09439_),
    .Y(_09446_));
 sky130_fd_sc_hd__nand3_4 _32001_ (.A(_09444_),
    .B(_09445_),
    .C(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__nor2_4 _32002_ (.A(_08986_),
    .B(_08981_),
    .Y(_09448_));
 sky130_fd_sc_hd__o2bb2ai_4 _32003_ (.A1_N(_09442_),
    .A2_N(_09447_),
    .B1(_08980_),
    .B2(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nor2_2 _32004_ (.A(_08980_),
    .B(_09448_),
    .Y(_09450_));
 sky130_fd_sc_hd__nand3_4 _32005_ (.A(_09447_),
    .B(_09442_),
    .C(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__nand2_1 _32006_ (.A(_09120_),
    .B(_09130_),
    .Y(_09452_));
 sky130_fd_sc_hd__nand2_4 _32007_ (.A(_09452_),
    .B(_09115_),
    .Y(_09453_));
 sky130_fd_sc_hd__a21oi_4 _32008_ (.A1(_09449_),
    .A2(_09451_),
    .B1(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__and3_1 _32009_ (.A(_09437_),
    .B(_09441_),
    .C(_09440_),
    .X(_09455_));
 sky130_fd_sc_hd__nand2_1 _32010_ (.A(_09447_),
    .B(_09450_),
    .Y(_09456_));
 sky130_fd_sc_hd__o211a_1 _32011_ (.A1(_09455_),
    .A2(_09456_),
    .B1(_09449_),
    .C1(_09453_),
    .X(_09457_));
 sky130_vsdinv _32012_ (.A(_08990_),
    .Y(_09458_));
 sky130_fd_sc_hd__and2_2 _32013_ (.A(_08995_),
    .B(_08998_),
    .X(_09459_));
 sky130_fd_sc_hd__nor2_4 _32014_ (.A(_09458_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__o21ai_2 _32015_ (.A1(_09454_),
    .A2(_09457_),
    .B1(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__a21o_1 _32016_ (.A1(_09449_),
    .A2(_09451_),
    .B1(_09453_),
    .X(_09462_));
 sky130_fd_sc_hd__nand3_4 _32017_ (.A(_09453_),
    .B(_09449_),
    .C(_09451_),
    .Y(_09463_));
 sky130_fd_sc_hd__nand3b_4 _32018_ (.A_N(_09460_),
    .B(_09462_),
    .C(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__a21oi_2 _32019_ (.A1(_08997_),
    .A2(_08999_),
    .B1(_08979_),
    .Y(_09465_));
 sky130_fd_sc_hd__o21ai_4 _32020_ (.A1(_09011_),
    .A2(_09465_),
    .B1(_09000_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand3_4 _32021_ (.A(_09461_),
    .B(_09464_),
    .C(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__o22ai_4 _32022_ (.A1(_09458_),
    .A2(_09459_),
    .B1(_09454_),
    .B2(_09457_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_1 _32023_ (.A(_09000_),
    .B(_09011_),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_2 _32024_ (.A(_09469_),
    .B(_09006_),
    .Y(_09470_));
 sky130_fd_sc_hd__nand3_2 _32025_ (.A(_09462_),
    .B(_09460_),
    .C(_09463_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand3_4 _32026_ (.A(_09468_),
    .B(_09470_),
    .C(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__nand2_1 _32027_ (.A(_09467_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__buf_6 _32028_ (.A(\pcpi_mul.rs1[27] ),
    .X(_09474_));
 sky130_fd_sc_hd__nand2_4 _32029_ (.A(_19937_),
    .B(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__clkbuf_4 _32030_ (.A(\pcpi_mul.rs1[23] ),
    .X(_09476_));
 sky130_fd_sc_hd__a22oi_4 _32031_ (.A1(_05228_),
    .A2(_08447_),
    .B1(_05367_),
    .B2(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__nor2_1 _32032_ (.A(_09475_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__nand2_2 _32033_ (.A(_06986_),
    .B(_08036_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2_2 _32034_ (.A(_06988_),
    .B(_08445_),
    .Y(_09480_));
 sky130_fd_sc_hd__or2_4 _32035_ (.A(_09479_),
    .B(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__nand2_2 _32036_ (.A(_09478_),
    .B(_09481_),
    .Y(_09482_));
 sky130_fd_sc_hd__nor2_4 _32037_ (.A(_09479_),
    .B(_09480_),
    .Y(_09483_));
 sky130_fd_sc_hd__o21ai_4 _32038_ (.A1(_09477_),
    .A2(_09483_),
    .B1(_09475_),
    .Y(_09484_));
 sky130_fd_sc_hd__o21ai_4 _32039_ (.A1(_09023_),
    .A2(_09026_),
    .B1(_09022_),
    .Y(_09485_));
 sky130_fd_sc_hd__a21oi_4 _32040_ (.A1(_09482_),
    .A2(_09484_),
    .B1(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__buf_4 _32041_ (.A(_09025_),
    .X(_09487_));
 sky130_fd_sc_hd__nand2_1 _32042_ (.A(_05240_),
    .B(_09038_),
    .Y(_09488_));
 sky130_fd_sc_hd__a21o_1 _32043_ (.A1(_05175_),
    .A2(_09487_),
    .B1(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__buf_6 _32044_ (.A(_09037_),
    .X(_09490_));
 sky130_fd_sc_hd__nand2_1 _32045_ (.A(_05242_),
    .B(_09025_),
    .Y(_09491_));
 sky130_fd_sc_hd__a21o_1 _32046_ (.A1(_05174_),
    .A2(_09490_),
    .B1(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__buf_6 _32047_ (.A(_20097_),
    .X(_09493_));
 sky130_fd_sc_hd__nand2_2 _32048_ (.A(_05830_),
    .B(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21oi_4 _32049_ (.A1(_09489_),
    .A2(_09492_),
    .B1(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__and3_1 _32050_ (.A(_09489_),
    .B(_09492_),
    .C(_09494_),
    .X(_09496_));
 sky130_fd_sc_hd__nor2_2 _32051_ (.A(_09495_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand3_4 _32052_ (.A(_09482_),
    .B(_09485_),
    .C(_09484_),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_1 _32053_ (.A(_09497_),
    .B(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__o21bai_2 _32054_ (.A1(_09477_),
    .A2(_09483_),
    .B1_N(_09475_),
    .Y(_09500_));
 sky130_vsdinv _32055_ (.A(_09477_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand3_2 _32056_ (.A(_09481_),
    .B(_09501_),
    .C(_09475_),
    .Y(_09502_));
 sky130_fd_sc_hd__o2111ai_4 _32057_ (.A1(_09023_),
    .A2(_09026_),
    .B1(_09022_),
    .C1(_09500_),
    .D1(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__nand2_1 _32058_ (.A(_09503_),
    .B(_09498_),
    .Y(_09504_));
 sky130_fd_sc_hd__a21o_1 _32059_ (.A1(_09489_),
    .A2(_09492_),
    .B1(_09494_),
    .X(_09505_));
 sky130_fd_sc_hd__nand3_1 _32060_ (.A(_09489_),
    .B(_09492_),
    .C(_09494_),
    .Y(_09506_));
 sky130_fd_sc_hd__nand2_2 _32061_ (.A(_09505_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__nand2_1 _32062_ (.A(_09504_),
    .B(_09507_),
    .Y(_09508_));
 sky130_fd_sc_hd__nand2_1 _32063_ (.A(_09062_),
    .B(_09036_),
    .Y(_09509_));
 sky130_fd_sc_hd__o211ai_4 _32064_ (.A1(_09486_),
    .A2(_09499_),
    .B1(_09508_),
    .C1(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__nand2_2 _32065_ (.A(_09504_),
    .B(_09497_),
    .Y(_09511_));
 sky130_fd_sc_hd__a21boi_4 _32066_ (.A1(_09049_),
    .A2(_09032_),
    .B1_N(_09036_),
    .Y(_09512_));
 sky130_fd_sc_hd__nand3_4 _32067_ (.A(_09503_),
    .B(_09507_),
    .C(_09498_),
    .Y(_09513_));
 sky130_fd_sc_hd__o21ba_1 _32068_ (.A1(_09039_),
    .A2(_09042_),
    .B1_N(_09046_),
    .X(_09514_));
 sky130_fd_sc_hd__a31oi_4 _32069_ (.A1(_09511_),
    .A2(_09512_),
    .A3(_09513_),
    .B1(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand3_2 _32070_ (.A(_09511_),
    .B(_09512_),
    .C(_09513_),
    .Y(_09516_));
 sky130_fd_sc_hd__a21boi_4 _32071_ (.A1(_09510_),
    .A2(_09516_),
    .B1_N(_09514_),
    .Y(_09517_));
 sky130_fd_sc_hd__a21oi_2 _32072_ (.A1(_09510_),
    .A2(_09515_),
    .B1(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__nand2_1 _32073_ (.A(_09473_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__and2_1 _32074_ (.A(_09515_),
    .B(_09510_),
    .X(_09520_));
 sky130_fd_sc_hd__o211ai_4 _32075_ (.A1(_09517_),
    .A2(_09520_),
    .B1(_09472_),
    .C1(_09467_),
    .Y(_09521_));
 sky130_fd_sc_hd__a21boi_4 _32076_ (.A1(_09142_),
    .A2(_09148_),
    .B1_N(_09146_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand3_4 _32077_ (.A(_09519_),
    .B(_09521_),
    .C(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__nand2_1 _32078_ (.A(_09142_),
    .B(_09148_),
    .Y(_09524_));
 sky130_fd_sc_hd__nand2_1 _32079_ (.A(_09524_),
    .B(_09146_),
    .Y(_09525_));
 sky130_fd_sc_hd__o2bb2ai_1 _32080_ (.A1_N(_09472_),
    .A2_N(_09467_),
    .B1(_09520_),
    .B2(_09517_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand3_1 _32081_ (.A(_09518_),
    .B(_09472_),
    .C(_09467_),
    .Y(_09527_));
 sky130_fd_sc_hd__nand3_2 _32082_ (.A(_09525_),
    .B(_09526_),
    .C(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__buf_2 _32083_ (.A(_09528_),
    .X(_09529_));
 sky130_vsdinv _32084_ (.A(_09014_),
    .Y(_09530_));
 sky130_fd_sc_hd__a21o_2 _32085_ (.A1(_09019_),
    .A2(_09066_),
    .B1(_09530_),
    .X(_09531_));
 sky130_fd_sc_hd__a21o_2 _32086_ (.A1(_09523_),
    .A2(_09529_),
    .B1(_09531_),
    .X(_09532_));
 sky130_fd_sc_hd__nand3_4 _32087_ (.A(_09523_),
    .B(_09529_),
    .C(_09531_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand3_2 _32088_ (.A(_09431_),
    .B(_09532_),
    .C(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__a21oi_4 _32089_ (.A1(_09523_),
    .A2(_09529_),
    .B1(_09531_),
    .Y(_09535_));
 sky130_fd_sc_hd__and2_1 _32090_ (.A(_09066_),
    .B(_09019_),
    .X(_09536_));
 sky130_fd_sc_hd__o211a_2 _32091_ (.A1(_09530_),
    .A2(_09536_),
    .B1(_09528_),
    .C1(_09523_),
    .X(_09537_));
 sky130_fd_sc_hd__o211ai_4 _32092_ (.A1(_09535_),
    .A2(_09537_),
    .B1(_09422_),
    .C1(_09430_),
    .Y(_09538_));
 sky130_fd_sc_hd__nand3_4 _32093_ (.A(_09267_),
    .B(_09534_),
    .C(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand3_1 _32094_ (.A(_09079_),
    .B(_09226_),
    .C(_09075_),
    .Y(_09540_));
 sky130_fd_sc_hd__nand2_2 _32095_ (.A(_09540_),
    .B(_09222_),
    .Y(_09541_));
 sky130_fd_sc_hd__o21ai_2 _32096_ (.A1(_09535_),
    .A2(_09537_),
    .B1(_09431_),
    .Y(_09542_));
 sky130_fd_sc_hd__nand2_2 _32097_ (.A(_09523_),
    .B(_09531_),
    .Y(_09543_));
 sky130_vsdinv _32098_ (.A(_09529_),
    .Y(_09544_));
 sky130_fd_sc_hd__o2111ai_4 _32099_ (.A1(_09543_),
    .A2(_09544_),
    .B1(_09430_),
    .C1(_09532_),
    .D1(_09422_),
    .Y(_09545_));
 sky130_fd_sc_hd__nand3_4 _32100_ (.A(_09541_),
    .B(_09542_),
    .C(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__a21oi_4 _32101_ (.A1(_09054_),
    .A2(_09056_),
    .B1(_09063_),
    .Y(_09547_));
 sky130_fd_sc_hd__a21oi_4 _32102_ (.A1(_09221_),
    .A2(_09068_),
    .B1(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__and3_2 _32103_ (.A(_09221_),
    .B(_09068_),
    .C(_09547_),
    .X(_09549_));
 sky130_fd_sc_hd__o2bb2ai_4 _32104_ (.A1_N(_09539_),
    .A2_N(_09546_),
    .B1(_09548_),
    .B2(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__nor2_4 _32105_ (.A(_09548_),
    .B(_09549_),
    .Y(_09551_));
 sky130_fd_sc_hd__nand3_4 _32106_ (.A(_09546_),
    .B(_09539_),
    .C(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__o21ai_4 _32107_ (.A1(_09235_),
    .A2(_09230_),
    .B1(_09239_),
    .Y(_09553_));
 sky130_fd_sc_hd__a21oi_4 _32108_ (.A1(_09550_),
    .A2(_09552_),
    .B1(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__a21oi_1 _32109_ (.A1(_09236_),
    .A2(_09237_),
    .B1(_09235_),
    .Y(_09555_));
 sky130_fd_sc_hd__o211a_1 _32110_ (.A1(_09233_),
    .A2(_09555_),
    .B1(_09552_),
    .C1(_09550_),
    .X(_09556_));
 sky130_fd_sc_hd__o21ai_1 _32111_ (.A1(_09554_),
    .A2(_09556_),
    .B1(_08970_),
    .Y(_09557_));
 sky130_fd_sc_hd__a21boi_2 _32112_ (.A1(_09248_),
    .A2(_08944_),
    .B1_N(_09244_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21o_1 _32113_ (.A1(_09550_),
    .A2(_09552_),
    .B1(_09553_),
    .X(_09559_));
 sky130_fd_sc_hd__nand3_4 _32114_ (.A(_09553_),
    .B(_09550_),
    .C(_09552_),
    .Y(_09560_));
 sky130_fd_sc_hd__nand3_2 _32115_ (.A(_09559_),
    .B(_08969_),
    .C(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__nand3_2 _32116_ (.A(_09557_),
    .B(_09558_),
    .C(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__o22ai_4 _32117_ (.A1(_08971_),
    .A2(_08968_),
    .B1(_09554_),
    .B2(_09556_),
    .Y(_09563_));
 sky130_fd_sc_hd__o21a_1 _32118_ (.A1(_09230_),
    .A2(_09233_),
    .B1(_09235_),
    .X(_09564_));
 sky130_fd_sc_hd__nand2_1 _32119_ (.A(_09240_),
    .B(_09243_),
    .Y(_09565_));
 sky130_fd_sc_hd__o2bb2ai_2 _32120_ (.A1_N(_08944_),
    .A2_N(_09248_),
    .B1(_09564_),
    .B2(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand3_2 _32121_ (.A(_09559_),
    .B(_08970_),
    .C(_09560_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand3_4 _32122_ (.A(_09563_),
    .B(_09566_),
    .C(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__and2_4 _32123_ (.A(_09562_),
    .B(_09568_),
    .X(_09569_));
 sky130_vsdinv _32124_ (.A(_09258_),
    .Y(_09570_));
 sky130_fd_sc_hd__o21ai_4 _32125_ (.A1(_09255_),
    .A2(_09266_),
    .B1(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__xor2_4 _32126_ (.A(_09569_),
    .B(_09571_),
    .X(_02646_));
 sky130_fd_sc_hd__o21ai_4 _32127_ (.A1(_08969_),
    .A2(_09554_),
    .B1(_09560_),
    .Y(_09572_));
 sky130_fd_sc_hd__nor2_2 _32128_ (.A(_09397_),
    .B(_09392_),
    .Y(_09573_));
 sky130_fd_sc_hd__nand2_2 _32129_ (.A(_07753_),
    .B(_06152_),
    .Y(_09574_));
 sky130_fd_sc_hd__nand2_2 _32130_ (.A(_06636_),
    .B(_20137_),
    .Y(_09575_));
 sky130_fd_sc_hd__nor2_4 _32131_ (.A(_09574_),
    .B(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__nand2_2 _32132_ (.A(_07893_),
    .B(_06441_),
    .Y(_09577_));
 sky130_vsdinv _32133_ (.A(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__nand2_2 _32134_ (.A(_09574_),
    .B(_09575_),
    .Y(_09579_));
 sky130_fd_sc_hd__nand3b_2 _32135_ (.A_N(_09576_),
    .B(_09578_),
    .C(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__a22oi_4 _32136_ (.A1(_07754_),
    .A2(_06153_),
    .B1(_06637_),
    .B2(_06309_),
    .Y(_09581_));
 sky130_fd_sc_hd__o21ai_2 _32137_ (.A1(_09581_),
    .A2(_09576_),
    .B1(_09577_),
    .Y(_09582_));
 sky130_fd_sc_hd__o22ai_4 _32138_ (.A1(_08242_),
    .A2(_09285_),
    .B1(_09287_),
    .B2(_09284_),
    .Y(_09583_));
 sky130_fd_sc_hd__nand3_4 _32139_ (.A(_09580_),
    .B(_09582_),
    .C(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__nand3b_2 _32140_ (.A_N(_09576_),
    .B(_09577_),
    .C(_09579_),
    .Y(_09585_));
 sky130_fd_sc_hd__a21oi_2 _32141_ (.A1(_09291_),
    .A2(_09293_),
    .B1(_09286_),
    .Y(_09586_));
 sky130_fd_sc_hd__o21ai_2 _32142_ (.A1(_09581_),
    .A2(_09576_),
    .B1(_09578_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand3_4 _32143_ (.A(_09585_),
    .B(_09586_),
    .C(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__nor2_8 _32144_ (.A(_09378_),
    .B(_09370_),
    .Y(_09589_));
 sky130_fd_sc_hd__o2bb2ai_4 _32145_ (.A1_N(_09584_),
    .A2_N(_09588_),
    .B1(_09369_),
    .B2(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__nor2_4 _32146_ (.A(_09369_),
    .B(_09589_),
    .Y(_09591_));
 sky130_fd_sc_hd__nand3_4 _32147_ (.A(_09588_),
    .B(_09584_),
    .C(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__nand2_4 _32148_ (.A(_09388_),
    .B(_09377_),
    .Y(_09593_));
 sky130_fd_sc_hd__a21oi_2 _32149_ (.A1(_09590_),
    .A2(_09592_),
    .B1(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__nand2_2 _32150_ (.A(_09588_),
    .B(_09591_),
    .Y(_09595_));
 sky130_vsdinv _32151_ (.A(_09584_),
    .Y(_09596_));
 sky130_fd_sc_hd__o211a_1 _32152_ (.A1(_09595_),
    .A2(_09596_),
    .B1(_09590_),
    .C1(_09593_),
    .X(_09597_));
 sky130_fd_sc_hd__a22oi_4 _32153_ (.A1(_19901_),
    .A2(_07702_),
    .B1(_19905_),
    .B2(_08042_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_4 _32154_ (.A(_06117_),
    .B(_20122_),
    .Y(_09599_));
 sky130_fd_sc_hd__nand2_4 _32155_ (.A(_06044_),
    .B(_07249_),
    .Y(_09600_));
 sky130_fd_sc_hd__nor2_8 _32156_ (.A(_09599_),
    .B(_09600_),
    .Y(_09601_));
 sky130_vsdinv _32157_ (.A(_07232_),
    .Y(_09602_));
 sky130_fd_sc_hd__nor2_4 _32158_ (.A(_05632_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__o21ai_1 _32159_ (.A1(_09598_),
    .A2(_09601_),
    .B1(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__nor2_1 _32160_ (.A(_09598_),
    .B(_09601_),
    .Y(_09605_));
 sky130_vsdinv _32161_ (.A(_09603_),
    .Y(_09606_));
 sky130_fd_sc_hd__nand2_1 _32162_ (.A(_09605_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__a21oi_4 _32163_ (.A1(_09341_),
    .A2(_09342_),
    .B1(_09346_),
    .Y(_09608_));
 sky130_fd_sc_hd__nand2_2 _32164_ (.A(_19892_),
    .B(_20132_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_2 _32165_ (.A(_06606_),
    .B(_06713_),
    .Y(_09610_));
 sky130_fd_sc_hd__or2_1 _32166_ (.A(_09609_),
    .B(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__nand2_1 _32167_ (.A(_07785_),
    .B(_20125_),
    .Y(_09612_));
 sky130_vsdinv _32168_ (.A(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__nand2_2 _32169_ (.A(_09609_),
    .B(_09610_),
    .Y(_09614_));
 sky130_fd_sc_hd__nand3_2 _32170_ (.A(_09611_),
    .B(_09613_),
    .C(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__a22oi_4 _32171_ (.A1(_06363_),
    .A2(_06715_),
    .B1(_06607_),
    .B2(_08002_),
    .Y(_09616_));
 sky130_fd_sc_hd__nor2_4 _32172_ (.A(_09609_),
    .B(_09610_),
    .Y(_09617_));
 sky130_fd_sc_hd__o21ai_2 _32173_ (.A1(_09616_),
    .A2(_09617_),
    .B1(_09612_),
    .Y(_09618_));
 sky130_fd_sc_hd__nand3b_4 _32174_ (.A_N(_09608_),
    .B(_09615_),
    .C(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__nand3_1 _32175_ (.A(_09611_),
    .B(_09612_),
    .C(_09614_),
    .Y(_09620_));
 sky130_fd_sc_hd__o21ai_1 _32176_ (.A1(_09616_),
    .A2(_09617_),
    .B1(_09613_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand3_2 _32177_ (.A(_09620_),
    .B(_09608_),
    .C(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__a22o_1 _32178_ (.A1(_09604_),
    .A2(_09607_),
    .B1(_09619_),
    .B2(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__nand2_1 _32179_ (.A(_09607_),
    .B(_09604_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand3b_1 _32180_ (.A_N(_09624_),
    .B(_09619_),
    .C(_09622_),
    .Y(_09625_));
 sky130_fd_sc_hd__nand2_2 _32181_ (.A(_09623_),
    .B(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__o21bai_4 _32182_ (.A1(_09594_),
    .A2(_09597_),
    .B1_N(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__a21o_1 _32183_ (.A1(_09590_),
    .A2(_09592_),
    .B1(_09593_),
    .X(_09628_));
 sky130_fd_sc_hd__nand3_4 _32184_ (.A(_09593_),
    .B(_09590_),
    .C(_09592_),
    .Y(_09629_));
 sky130_fd_sc_hd__nand3_4 _32185_ (.A(_09628_),
    .B(_09629_),
    .C(_09626_),
    .Y(_09630_));
 sky130_fd_sc_hd__o21ai_4 _32186_ (.A1(_09329_),
    .A2(_09297_),
    .B1(_09298_),
    .Y(_09631_));
 sky130_fd_sc_hd__a21oi_4 _32187_ (.A1(_09627_),
    .A2(_09630_),
    .B1(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__nor2_1 _32188_ (.A(_09329_),
    .B(_09297_),
    .Y(_09633_));
 sky130_fd_sc_hd__o211a_2 _32189_ (.A1(_09328_),
    .A2(_09633_),
    .B1(_09630_),
    .C1(_09627_),
    .X(_09634_));
 sky130_fd_sc_hd__o22ai_2 _32190_ (.A1(_09390_),
    .A2(_09573_),
    .B1(_09632_),
    .B2(_09634_),
    .Y(_09635_));
 sky130_fd_sc_hd__nand2_2 _32191_ (.A(_09627_),
    .B(_09630_),
    .Y(_09636_));
 sky130_vsdinv _32192_ (.A(_09631_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand2_2 _32193_ (.A(_09636_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__nand3_2 _32194_ (.A(_09627_),
    .B(_09630_),
    .C(_09631_),
    .Y(_09639_));
 sky130_fd_sc_hd__a21oi_4 _32195_ (.A1(_09394_),
    .A2(_09397_),
    .B1(_09392_),
    .Y(_09640_));
 sky130_vsdinv _32196_ (.A(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__nand3_1 _32197_ (.A(_09638_),
    .B(_09639_),
    .C(_09641_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand2_1 _32198_ (.A(_09635_),
    .B(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__a22oi_4 _32199_ (.A1(_08589_),
    .A2(_05218_),
    .B1(_08575_),
    .B2(_07417_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand3_4 _32200_ (.A(_19857_),
    .B(_08761_),
    .C(_05285_),
    .Y(_09645_));
 sky130_fd_sc_hd__nor2_8 _32201_ (.A(_05295_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand2_4 _32202_ (.A(\pcpi_mul.rs2[21] ),
    .B(_05372_),
    .Y(_09647_));
 sky130_vsdinv _32203_ (.A(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__o21ai_2 _32204_ (.A1(_09644_),
    .A2(_09646_),
    .B1(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21oi_2 _32205_ (.A1(_09277_),
    .A2(_09276_),
    .B1(_09271_),
    .Y(_09650_));
 sky130_fd_sc_hd__a22o_1 _32206_ (.A1(_08589_),
    .A2(_05392_),
    .B1(_08575_),
    .B2(_07417_),
    .X(_09651_));
 sky130_fd_sc_hd__o211ai_2 _32207_ (.A1(_05580_),
    .A2(_09645_),
    .B1(_09647_),
    .C1(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__nand3_4 _32208_ (.A(_09649_),
    .B(_09650_),
    .C(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__nand2_1 _32209_ (.A(_09651_),
    .B(_09648_),
    .Y(_09654_));
 sky130_fd_sc_hd__o22ai_4 _32210_ (.A1(_09275_),
    .A2(_09270_),
    .B1(_09272_),
    .B2(_09268_),
    .Y(_09655_));
 sky130_fd_sc_hd__o21ai_2 _32211_ (.A1(_09644_),
    .A2(_09646_),
    .B1(_09647_),
    .Y(_09656_));
 sky130_fd_sc_hd__o211ai_4 _32212_ (.A1(_09646_),
    .A2(_09654_),
    .B1(_09655_),
    .C1(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand2_1 _32213_ (.A(_19869_),
    .B(_06475_),
    .Y(_09658_));
 sky130_fd_sc_hd__nand3b_4 _32214_ (.A_N(_09658_),
    .B(_08248_),
    .C(_06289_),
    .Y(_09659_));
 sky130_fd_sc_hd__a22o_2 _32215_ (.A1(_08326_),
    .A2(_05698_),
    .B1(_19873_),
    .B2(_05699_),
    .X(_09660_));
 sky130_fd_sc_hd__nand2_2 _32216_ (.A(_19876_),
    .B(_20145_),
    .Y(_09661_));
 sky130_vsdinv _32217_ (.A(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__a21oi_2 _32218_ (.A1(_09659_),
    .A2(_09660_),
    .B1(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__and3_1 _32219_ (.A(_09659_),
    .B(_09662_),
    .C(_09660_),
    .X(_09664_));
 sky130_fd_sc_hd__o2bb2ai_4 _32220_ (.A1_N(_09653_),
    .A2_N(_09657_),
    .B1(_09663_),
    .B2(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__a22oi_4 _32221_ (.A1(_07482_),
    .A2(_05831_),
    .B1(_08248_),
    .B2(_20149_),
    .Y(_09666_));
 sky130_fd_sc_hd__and4_1 _32222_ (.A(_08779_),
    .B(_08598_),
    .C(_06480_),
    .D(_05454_),
    .X(_09667_));
 sky130_fd_sc_hd__o21ai_1 _32223_ (.A1(_09666_),
    .A2(_09667_),
    .B1(_09662_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand3_1 _32224_ (.A(_09659_),
    .B(_09661_),
    .C(_09660_),
    .Y(_09669_));
 sky130_fd_sc_hd__nand2_2 _32225_ (.A(_09668_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand3_4 _32226_ (.A(_09657_),
    .B(_09653_),
    .C(_09670_),
    .Y(_09671_));
 sky130_fd_sc_hd__nand2_1 _32227_ (.A(_09312_),
    .B(_09314_),
    .Y(_09672_));
 sky130_fd_sc_hd__nor2_4 _32228_ (.A(_09304_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__a21oi_4 _32229_ (.A1(_09665_),
    .A2(_09671_),
    .B1(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__and3_2 _32230_ (.A(_09665_),
    .B(_09673_),
    .C(_09671_),
    .X(_09675_));
 sky130_fd_sc_hd__nand2_4 _32231_ (.A(_09296_),
    .B(_09279_),
    .Y(_09676_));
 sky130_vsdinv _32232_ (.A(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__o21ai_4 _32233_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__nand2_2 _32234_ (.A(_19846_),
    .B(_05125_),
    .Y(_09679_));
 sky130_fd_sc_hd__nand2_2 _32235_ (.A(_08799_),
    .B(_20167_),
    .Y(_09680_));
 sky130_fd_sc_hd__nor2_4 _32236_ (.A(_09679_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__and2_1 _32237_ (.A(_09679_),
    .B(_09680_),
    .X(_09682_));
 sky130_fd_sc_hd__nand2_2 _32238_ (.A(\pcpi_mul.rs2[24] ),
    .B(_05251_),
    .Y(_09683_));
 sky130_fd_sc_hd__o21ai_2 _32239_ (.A1(_09681_),
    .A2(_09682_),
    .B1(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__or2_2 _32240_ (.A(_09679_),
    .B(_09680_),
    .X(_09685_));
 sky130_fd_sc_hd__nand2_2 _32241_ (.A(_09679_),
    .B(_09680_),
    .Y(_09686_));
 sky130_vsdinv _32242_ (.A(_09683_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand3_2 _32243_ (.A(_09685_),
    .B(_09686_),
    .C(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__a31o_1 _32244_ (.A1(_09308_),
    .A2(_08802_),
    .A3(_06614_),
    .B1(_09307_),
    .X(_09689_));
 sky130_fd_sc_hd__nand3_4 _32245_ (.A(_09684_),
    .B(_09688_),
    .C(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__o21ai_2 _32246_ (.A1(_09681_),
    .A2(_09682_),
    .B1(_09687_),
    .Y(_09691_));
 sky130_fd_sc_hd__nand3_2 _32247_ (.A(_09685_),
    .B(_09686_),
    .C(_09683_),
    .Y(_09692_));
 sky130_fd_sc_hd__a21oi_2 _32248_ (.A1(_09310_),
    .A2(_09308_),
    .B1(_09307_),
    .Y(_09693_));
 sky130_fd_sc_hd__nand3_4 _32249_ (.A(_09691_),
    .B(_09692_),
    .C(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__nand2_2 _32250_ (.A(_19839_),
    .B(_20176_),
    .Y(_09695_));
 sky130_fd_sc_hd__buf_4 _32251_ (.A(\pcpi_mul.rs2[27] ),
    .X(_09696_));
 sky130_fd_sc_hd__nand2_2 _32252_ (.A(_09696_),
    .B(_20173_),
    .Y(_09697_));
 sky130_fd_sc_hd__nor2_8 _32253_ (.A(_09695_),
    .B(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__and2_2 _32254_ (.A(_09695_),
    .B(_09697_),
    .X(_09699_));
 sky130_fd_sc_hd__nor2_4 _32255_ (.A(_09698_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__a21oi_2 _32256_ (.A1(_09690_),
    .A2(_09694_),
    .B1(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__nor2_1 _32257_ (.A(_09325_),
    .B(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__nand3_4 _32258_ (.A(_09690_),
    .B(_09694_),
    .C(_09700_),
    .Y(_09703_));
 sky130_fd_sc_hd__o2bb2ai_1 _32259_ (.A1_N(_09694_),
    .A2_N(_09690_),
    .B1(_09698_),
    .B2(_09699_),
    .Y(_09704_));
 sky130_fd_sc_hd__a21boi_1 _32260_ (.A1(_09704_),
    .A2(_09703_),
    .B1_N(_09325_),
    .Y(_09705_));
 sky130_fd_sc_hd__a21oi_2 _32261_ (.A1(_09702_),
    .A2(_09703_),
    .B1(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__nand2_1 _32262_ (.A(_09665_),
    .B(_09671_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand2_2 _32263_ (.A(_09707_),
    .B(_09315_),
    .Y(_09708_));
 sky130_fd_sc_hd__nand3_4 _32264_ (.A(_09665_),
    .B(_09673_),
    .C(_09671_),
    .Y(_09709_));
 sky130_fd_sc_hd__nand3_4 _32265_ (.A(_09708_),
    .B(_09676_),
    .C(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__nand3_4 _32266_ (.A(_09678_),
    .B(_09706_),
    .C(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__o21ai_2 _32267_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09676_),
    .Y(_09712_));
 sky130_fd_sc_hd__nand2_1 _32268_ (.A(_09702_),
    .B(_09703_),
    .Y(_09713_));
 sky130_vsdinv _32269_ (.A(_09703_),
    .Y(_09714_));
 sky130_fd_sc_hd__o21ai_2 _32270_ (.A1(_09701_),
    .A2(_09714_),
    .B1(_09325_),
    .Y(_09715_));
 sky130_fd_sc_hd__nand2_1 _32271_ (.A(_09713_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__nand3_2 _32272_ (.A(_09708_),
    .B(_09677_),
    .C(_09709_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand3_4 _32273_ (.A(_09712_),
    .B(_09716_),
    .C(_09717_),
    .Y(_09718_));
 sky130_fd_sc_hd__o2bb2ai_1 _32274_ (.A1_N(_09711_),
    .A2_N(_09718_),
    .B1(_09301_),
    .B2(_09335_),
    .Y(_09719_));
 sky130_fd_sc_hd__nand3b_4 _32275_ (.A_N(_09333_),
    .B(_09711_),
    .C(_09718_),
    .Y(_09720_));
 sky130_fd_sc_hd__nand2_1 _32276_ (.A(_09719_),
    .B(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__nand2_2 _32277_ (.A(_09643_),
    .B(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__o21ai_4 _32278_ (.A1(_09334_),
    .A2(_09417_),
    .B1(_09420_),
    .Y(_09723_));
 sky130_vsdinv _32279_ (.A(_09711_),
    .Y(_09724_));
 sky130_fd_sc_hd__nor2_2 _32280_ (.A(_09326_),
    .B(_09303_),
    .Y(_09725_));
 sky130_fd_sc_hd__nand3_4 _32281_ (.A(_09718_),
    .B(_09725_),
    .C(_09331_),
    .Y(_09726_));
 sky130_fd_sc_hd__clkbuf_4 _32282_ (.A(_09719_),
    .X(_09727_));
 sky130_fd_sc_hd__clkbuf_4 _32283_ (.A(_09642_),
    .X(_09728_));
 sky130_fd_sc_hd__clkbuf_4 _32284_ (.A(_09635_),
    .X(_09729_));
 sky130_fd_sc_hd__o2111ai_4 _32285_ (.A1(_09724_),
    .A2(_09726_),
    .B1(_09727_),
    .C1(_09728_),
    .D1(_09729_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand3_2 _32286_ (.A(_09722_),
    .B(_09723_),
    .C(_09730_),
    .Y(_09731_));
 sky130_vsdinv _32287_ (.A(\pcpi_mul.rs1[21] ),
    .Y(_09732_));
 sky130_fd_sc_hd__buf_6 _32288_ (.A(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__nand3_4 _32289_ (.A(_05502_),
    .B(_05413_),
    .C(_20110_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_2 _32290_ (.A(_05506_),
    .B(_20104_),
    .Y(_09735_));
 sky130_fd_sc_hd__a22oi_4 _32291_ (.A1(_05502_),
    .A2(_07548_),
    .B1(_05499_),
    .B2(_08057_),
    .Y(_09736_));
 sky130_fd_sc_hd__nor2_4 _32292_ (.A(_09735_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__o21ai_2 _32293_ (.A1(_09733_),
    .A2(_09734_),
    .B1(_09737_),
    .Y(_09738_));
 sky130_fd_sc_hd__a21o_1 _32294_ (.A1(_09361_),
    .A2(_09357_),
    .B1(_09360_),
    .X(_09739_));
 sky130_fd_sc_hd__nor2_4 _32295_ (.A(_09732_),
    .B(_09734_),
    .Y(_09740_));
 sky130_fd_sc_hd__o21ai_2 _32296_ (.A1(_09736_),
    .A2(_09740_),
    .B1(_09735_),
    .Y(_09741_));
 sky130_fd_sc_hd__nand3_4 _32297_ (.A(_09738_),
    .B(_09739_),
    .C(_09741_),
    .Y(_09742_));
 sky130_vsdinv _32298_ (.A(_09736_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand3b_2 _32299_ (.A_N(_09740_),
    .B(_09743_),
    .C(_09735_),
    .Y(_09744_));
 sky130_fd_sc_hd__a21oi_4 _32300_ (.A1(_09361_),
    .A2(_09357_),
    .B1(_09360_),
    .Y(_09745_));
 sky130_fd_sc_hd__o21bai_2 _32301_ (.A1(_09736_),
    .A2(_09740_),
    .B1_N(_09735_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand3_4 _32302_ (.A(_09744_),
    .B(_09745_),
    .C(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__nor2_4 _32303_ (.A(_09438_),
    .B(_09435_),
    .Y(_09748_));
 sky130_fd_sc_hd__o2bb2ai_4 _32304_ (.A1_N(_09742_),
    .A2_N(_09747_),
    .B1(_09432_),
    .B2(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__nor2_4 _32305_ (.A(_09432_),
    .B(_09748_),
    .Y(_09750_));
 sky130_fd_sc_hd__nand3_4 _32306_ (.A(_09747_),
    .B(_09742_),
    .C(_09750_),
    .Y(_09751_));
 sky130_vsdinv _32307_ (.A(_09347_),
    .Y(_09752_));
 sky130_fd_sc_hd__nand2_1 _32308_ (.A(_09343_),
    .B(_09344_),
    .Y(_09753_));
 sky130_fd_sc_hd__o2bb2ai_4 _32309_ (.A1_N(_09363_),
    .A2_N(_09352_),
    .B1(_09752_),
    .B2(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__a21oi_4 _32310_ (.A1(_09749_),
    .A2(_09751_),
    .B1(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_1 _32311_ (.A(_09747_),
    .B(_09750_),
    .Y(_09756_));
 sky130_vsdinv _32312_ (.A(_09742_),
    .Y(_09757_));
 sky130_fd_sc_hd__o211a_1 _32313_ (.A1(_09756_),
    .A2(_09757_),
    .B1(_09754_),
    .C1(_09749_),
    .X(_09758_));
 sky130_vsdinv _32314_ (.A(_09451_),
    .Y(_09759_));
 sky130_fd_sc_hd__nor2_2 _32315_ (.A(_09455_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__clkbuf_2 _32316_ (.A(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__o21bai_2 _32317_ (.A1(_09755_),
    .A2(_09758_),
    .B1_N(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__o21a_1 _32318_ (.A1(_09460_),
    .A2(_09454_),
    .B1(_09463_),
    .X(_09763_));
 sky130_vsdinv _32319_ (.A(_09754_),
    .Y(_09764_));
 sky130_fd_sc_hd__nand2_1 _32320_ (.A(_09749_),
    .B(_09751_),
    .Y(_09765_));
 sky130_fd_sc_hd__nand2_2 _32321_ (.A(_09764_),
    .B(_09765_),
    .Y(_09766_));
 sky130_fd_sc_hd__nand3_4 _32322_ (.A(_09749_),
    .B(_09754_),
    .C(_09751_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand3_2 _32323_ (.A(_09766_),
    .B(_09767_),
    .C(_09761_),
    .Y(_09768_));
 sky130_fd_sc_hd__nand3_4 _32324_ (.A(_09762_),
    .B(_09763_),
    .C(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__o21ai_2 _32325_ (.A1(_09755_),
    .A2(_09758_),
    .B1(_09761_),
    .Y(_09770_));
 sky130_fd_sc_hd__nand3b_2 _32326_ (.A_N(_09760_),
    .B(_09766_),
    .C(_09767_),
    .Y(_09771_));
 sky130_fd_sc_hd__o21ai_2 _32327_ (.A1(_09460_),
    .A2(_09454_),
    .B1(_09463_),
    .Y(_09772_));
 sky130_fd_sc_hd__nand3_4 _32328_ (.A(_09770_),
    .B(_09771_),
    .C(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__o21ai_2 _32329_ (.A1(_09507_),
    .A2(_09486_),
    .B1(_09498_),
    .Y(_09774_));
 sky130_vsdinv _32330_ (.A(\pcpi_mul.rs1[28] ),
    .Y(_09775_));
 sky130_fd_sc_hd__nand3_4 _32331_ (.A(_05311_),
    .B(_05377_),
    .C(_08445_),
    .Y(_09776_));
 sky130_fd_sc_hd__a22o_2 _32332_ (.A1(_05450_),
    .A2(_09476_),
    .B1(_05367_),
    .B2(_20096_),
    .X(_09777_));
 sky130_fd_sc_hd__o21ai_2 _32333_ (.A1(_08435_),
    .A2(_09776_),
    .B1(_09777_),
    .Y(_09778_));
 sky130_fd_sc_hd__o21ai_4 _32334_ (.A1(_04837_),
    .A2(_09775_),
    .B1(_09778_),
    .Y(_09779_));
 sky130_fd_sc_hd__nor2_1 _32335_ (.A(_08435_),
    .B(_09776_),
    .Y(_09780_));
 sky130_fd_sc_hd__nor2_2 _32336_ (.A(_04836_),
    .B(_09775_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand3b_4 _32337_ (.A_N(_09780_),
    .B(_09777_),
    .C(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__o21ai_4 _32338_ (.A1(_09475_),
    .A2(_09477_),
    .B1(_09481_),
    .Y(_09783_));
 sky130_fd_sc_hd__a21oi_4 _32339_ (.A1(_09779_),
    .A2(_09782_),
    .B1(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__nand3_4 _32340_ (.A(_09779_),
    .B(_09783_),
    .C(_09782_),
    .Y(_09785_));
 sky130_vsdinv _32341_ (.A(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__buf_6 _32342_ (.A(_20085_),
    .X(_09787_));
 sky130_fd_sc_hd__nand2_2 _32343_ (.A(_06314_),
    .B(_20090_),
    .Y(_09788_));
 sky130_fd_sc_hd__a21o_1 _32344_ (.A1(_05175_),
    .A2(_09787_),
    .B1(_09788_),
    .X(_09789_));
 sky130_fd_sc_hd__nand2_2 _32345_ (.A(_19934_),
    .B(_09474_),
    .Y(_09790_));
 sky130_fd_sc_hd__a21o_1 _32346_ (.A1(_05174_),
    .A2(_09487_),
    .B1(_09790_),
    .X(_09791_));
 sky130_fd_sc_hd__nand2_2 _32347_ (.A(_19928_),
    .B(_20094_),
    .Y(_09792_));
 sky130_fd_sc_hd__a21o_1 _32348_ (.A1(_09789_),
    .A2(_09791_),
    .B1(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__nand3_2 _32349_ (.A(_09789_),
    .B(_09791_),
    .C(_09792_),
    .Y(_09794_));
 sky130_fd_sc_hd__and2_1 _32350_ (.A(_09793_),
    .B(_09794_),
    .X(_09795_));
 sky130_fd_sc_hd__o21ai_2 _32351_ (.A1(_09784_),
    .A2(_09786_),
    .B1(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__a21o_1 _32352_ (.A1(_09779_),
    .A2(_09782_),
    .B1(_09783_),
    .X(_09797_));
 sky130_fd_sc_hd__nand2_2 _32353_ (.A(_09793_),
    .B(_09794_),
    .Y(_09798_));
 sky130_fd_sc_hd__nand3_2 _32354_ (.A(_09797_),
    .B(_09798_),
    .C(_09785_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand3b_4 _32355_ (.A_N(_09774_),
    .B(_09796_),
    .C(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_1 _32356_ (.A(_09795_),
    .B(_09797_),
    .Y(_09801_));
 sky130_fd_sc_hd__o21ai_2 _32357_ (.A1(_09784_),
    .A2(_09786_),
    .B1(_09798_),
    .Y(_09802_));
 sky130_fd_sc_hd__o211ai_4 _32358_ (.A1(_09786_),
    .A2(_09801_),
    .B1(_09774_),
    .C1(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__nor2_2 _32359_ (.A(_09488_),
    .B(_09491_),
    .Y(_09804_));
 sky130_fd_sc_hd__or2_4 _32360_ (.A(_09804_),
    .B(_09495_),
    .X(_09805_));
 sky130_fd_sc_hd__and3_1 _32361_ (.A(_09800_),
    .B(_09803_),
    .C(_09805_),
    .X(_09806_));
 sky130_fd_sc_hd__a21oi_4 _32362_ (.A1(_09800_),
    .A2(_09803_),
    .B1(_09805_),
    .Y(_09807_));
 sky130_fd_sc_hd__o2bb2ai_4 _32363_ (.A1_N(_09769_),
    .A2_N(_09773_),
    .B1(_09806_),
    .B2(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__o2bb2ai_1 _32364_ (.A1_N(_09803_),
    .A2_N(_09800_),
    .B1(_09804_),
    .B2(_09495_),
    .Y(_09809_));
 sky130_fd_sc_hd__nand3b_1 _32365_ (.A_N(_09805_),
    .B(_09800_),
    .C(_09803_),
    .Y(_09810_));
 sky130_fd_sc_hd__nand2_2 _32366_ (.A(_09809_),
    .B(_09810_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand3_4 _32367_ (.A(_09811_),
    .B(_09769_),
    .C(_09773_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2_2 _32368_ (.A(_09427_),
    .B(_09401_),
    .Y(_09813_));
 sky130_fd_sc_hd__a21o_1 _32369_ (.A1(_09808_),
    .A2(_09812_),
    .B1(_09813_),
    .X(_09814_));
 sky130_fd_sc_hd__nand3_4 _32370_ (.A(_09808_),
    .B(_09813_),
    .C(_09812_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_1 _32371_ (.A(_09518_),
    .B(_09472_),
    .Y(_09816_));
 sky130_fd_sc_hd__nand2_2 _32372_ (.A(_09816_),
    .B(_09467_),
    .Y(_09817_));
 sky130_fd_sc_hd__nand3_4 _32373_ (.A(_09814_),
    .B(_09815_),
    .C(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__and2_1 _32374_ (.A(_09731_),
    .B(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__nand2_1 _32375_ (.A(_09814_),
    .B(_09815_),
    .Y(_09820_));
 sky130_vsdinv _32376_ (.A(_09817_),
    .Y(_09821_));
 sky130_fd_sc_hd__nand2_1 _32377_ (.A(_09722_),
    .B(_09730_),
    .Y(_09822_));
 sky130_vsdinv _32378_ (.A(_09723_),
    .Y(_09823_));
 sky130_fd_sc_hd__a22oi_4 _32379_ (.A1(_09820_),
    .A2(_09821_),
    .B1(_09822_),
    .B2(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_1 _32380_ (.A(_09819_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__a21oi_4 _32381_ (.A1(_09722_),
    .A2(_09730_),
    .B1(_09723_),
    .Y(_09826_));
 sky130_fd_sc_hd__nand3_1 _32382_ (.A(_09728_),
    .B(_09727_),
    .C(_09720_),
    .Y(_09827_));
 sky130_vsdinv _32383_ (.A(_09729_),
    .Y(_09828_));
 sky130_fd_sc_hd__o211a_2 _32384_ (.A1(_09827_),
    .A2(_09828_),
    .B1(_09723_),
    .C1(_09722_),
    .X(_09829_));
 sky130_fd_sc_hd__a21oi_2 _32385_ (.A1(_09808_),
    .A2(_09812_),
    .B1(_09813_),
    .Y(_09830_));
 sky130_fd_sc_hd__o211a_1 _32386_ (.A1(_09426_),
    .A2(_09407_),
    .B1(_09812_),
    .C1(_09808_),
    .X(_09831_));
 sky130_fd_sc_hd__o21ai_4 _32387_ (.A1(_09830_),
    .A2(_09831_),
    .B1(_09821_),
    .Y(_09832_));
 sky130_fd_sc_hd__nand2_4 _32388_ (.A(_09832_),
    .B(_09818_),
    .Y(_09833_));
 sky130_fd_sc_hd__o21ai_4 _32389_ (.A1(_09826_),
    .A2(_09829_),
    .B1(_09833_),
    .Y(_09834_));
 sky130_fd_sc_hd__and3_1 _32390_ (.A(_09425_),
    .B(_09428_),
    .C(_09429_),
    .X(_09835_));
 sky130_fd_sc_hd__a31o_1 _32391_ (.A1(_09532_),
    .A2(_09533_),
    .A3(_09422_),
    .B1(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__nand3_4 _32392_ (.A(_09825_),
    .B(_09834_),
    .C(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__a22oi_4 _32393_ (.A1(_09727_),
    .A2(_09720_),
    .B1(_09729_),
    .B2(_09728_),
    .Y(_09838_));
 sky130_fd_sc_hd__o2111a_1 _32394_ (.A1(_09724_),
    .A2(_09726_),
    .B1(_09727_),
    .C1(_09728_),
    .D1(_09729_),
    .X(_09839_));
 sky130_fd_sc_hd__o21bai_4 _32395_ (.A1(_09838_),
    .A2(_09839_),
    .B1_N(_09723_),
    .Y(_09840_));
 sky130_fd_sc_hd__a21o_1 _32396_ (.A1(_09840_),
    .A2(_09731_),
    .B1(_09833_),
    .X(_09841_));
 sky130_fd_sc_hd__a31oi_4 _32397_ (.A1(_09533_),
    .A2(_09532_),
    .A3(_09422_),
    .B1(_09835_),
    .Y(_09842_));
 sky130_fd_sc_hd__nand3_2 _32398_ (.A(_09833_),
    .B(_09840_),
    .C(_09731_),
    .Y(_09843_));
 sky130_fd_sc_hd__nand3_4 _32399_ (.A(_09841_),
    .B(_09842_),
    .C(_09843_),
    .Y(_09844_));
 sky130_vsdinv _32400_ (.A(_09515_),
    .Y(_09845_));
 sky130_fd_sc_hd__nand2_1 _32401_ (.A(_09845_),
    .B(_09510_),
    .Y(_09846_));
 sky130_vsdinv _32402_ (.A(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__nor2_4 _32403_ (.A(_09544_),
    .B(_09537_),
    .Y(_09848_));
 sky130_fd_sc_hd__nor2_8 _32404_ (.A(_09847_),
    .B(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__and3_1 _32405_ (.A(_09543_),
    .B(_09529_),
    .C(_09847_),
    .X(_09850_));
 sky130_fd_sc_hd__o2bb2ai_1 _32406_ (.A1_N(_09837_),
    .A2_N(_09844_),
    .B1(_09849_),
    .B2(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__nor2_4 _32407_ (.A(_09850_),
    .B(_09849_),
    .Y(_09852_));
 sky130_fd_sc_hd__nand3_1 _32408_ (.A(_09844_),
    .B(_09837_),
    .C(_09852_),
    .Y(_09853_));
 sky130_fd_sc_hd__nand2_1 _32409_ (.A(_09552_),
    .B(_09546_),
    .Y(_09854_));
 sky130_fd_sc_hd__nand3_2 _32410_ (.A(_09851_),
    .B(_09853_),
    .C(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__buf_2 _32411_ (.A(_09855_),
    .X(_09856_));
 sky130_fd_sc_hd__nor2_1 _32412_ (.A(_09846_),
    .B(_09848_),
    .Y(_09857_));
 sky130_fd_sc_hd__and3_1 _32413_ (.A(_09543_),
    .B(_09529_),
    .C(_09846_),
    .X(_09858_));
 sky130_fd_sc_hd__o2bb2ai_1 _32414_ (.A1_N(_09837_),
    .A2_N(_09844_),
    .B1(_09857_),
    .B2(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__a21boi_2 _32415_ (.A1(_09551_),
    .A2(_09539_),
    .B1_N(_09546_),
    .Y(_09860_));
 sky130_fd_sc_hd__nand3b_2 _32416_ (.A_N(_09852_),
    .B(_09844_),
    .C(_09837_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand3_2 _32417_ (.A(_09859_),
    .B(_09860_),
    .C(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__buf_2 _32418_ (.A(_09548_),
    .X(_09863_));
 sky130_fd_sc_hd__a21bo_1 _32419_ (.A1(_09856_),
    .A2(_09862_),
    .B1_N(_09863_),
    .X(_09864_));
 sky130_fd_sc_hd__clkbuf_4 _32420_ (.A(_09862_),
    .X(_09865_));
 sky130_fd_sc_hd__nand3b_2 _32421_ (.A_N(_09548_),
    .B(_09856_),
    .C(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__nand3b_4 _32422_ (.A_N(_09572_),
    .B(_09864_),
    .C(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__a21o_1 _32423_ (.A1(_09856_),
    .A2(_09865_),
    .B1(_09863_),
    .X(_09868_));
 sky130_fd_sc_hd__nand3_2 _32424_ (.A(_09856_),
    .B(_09865_),
    .C(_09863_),
    .Y(_09869_));
 sky130_fd_sc_hd__nand3_2 _32425_ (.A(_09868_),
    .B(_09572_),
    .C(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__nand2_1 _32426_ (.A(_09867_),
    .B(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__nand3_4 _32427_ (.A(_09264_),
    .B(_09569_),
    .C(_09259_),
    .Y(_09872_));
 sky130_fd_sc_hd__nand3_2 _32428_ (.A(_09260_),
    .B(_09569_),
    .C(_09259_),
    .Y(_09873_));
 sky130_fd_sc_hd__nand2_1 _32429_ (.A(_09258_),
    .B(_09562_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand3_4 _32430_ (.A(_09873_),
    .B(_09568_),
    .C(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__o21bai_4 _32431_ (.A1(_09872_),
    .A2(_08682_),
    .B1_N(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__xnor2_2 _32432_ (.A(_09871_),
    .B(_09876_),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _32433_ (.A(_09844_),
    .B(_09852_),
    .Y(_09877_));
 sky130_fd_sc_hd__nand2_2 _32434_ (.A(_09877_),
    .B(_09837_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand2_2 _32435_ (.A(_09639_),
    .B(_09640_),
    .Y(_09879_));
 sky130_fd_sc_hd__clkbuf_8 _32436_ (.A(_08888_),
    .X(_09880_));
 sky130_fd_sc_hd__nand2_2 _32437_ (.A(_05450_),
    .B(_20096_),
    .Y(_09881_));
 sky130_fd_sc_hd__nand2_2 _32438_ (.A(_05367_),
    .B(_09037_),
    .Y(_09882_));
 sky130_fd_sc_hd__or2_1 _32439_ (.A(_09881_),
    .B(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__nand2_2 _32440_ (.A(_05217_),
    .B(_20077_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand2_2 _32441_ (.A(_09881_),
    .B(_09882_),
    .Y(_09885_));
 sky130_fd_sc_hd__nand3_2 _32442_ (.A(_09883_),
    .B(_09884_),
    .C(_09885_),
    .Y(_09886_));
 sky130_fd_sc_hd__nor2_4 _32443_ (.A(_09881_),
    .B(_09882_),
    .Y(_09887_));
 sky130_fd_sc_hd__and2_1 _32444_ (.A(_09881_),
    .B(_09882_),
    .X(_09888_));
 sky130_vsdinv _32445_ (.A(_09884_),
    .Y(_09889_));
 sky130_fd_sc_hd__o21ai_2 _32446_ (.A1(_09887_),
    .A2(_09888_),
    .B1(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__o2111ai_4 _32447_ (.A1(_09880_),
    .A2(_09776_),
    .B1(_09782_),
    .C1(_09886_),
    .D1(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__a21o_1 _32448_ (.A1(_09781_),
    .A2(_09777_),
    .B1(_09780_),
    .X(_09892_));
 sky130_fd_sc_hd__o21ai_2 _32449_ (.A1(_09887_),
    .A2(_09888_),
    .B1(_09884_),
    .Y(_09893_));
 sky130_fd_sc_hd__nand3_2 _32450_ (.A(_09883_),
    .B(_09889_),
    .C(_09885_),
    .Y(_09894_));
 sky130_fd_sc_hd__nand3_4 _32451_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .Y(_09895_));
 sky130_fd_sc_hd__buf_6 _32452_ (.A(_20081_),
    .X(_09896_));
 sky130_fd_sc_hd__nand2_1 _32453_ (.A(_19931_),
    .B(_09474_),
    .Y(_09897_));
 sky130_fd_sc_hd__a21o_1 _32454_ (.A1(_05175_),
    .A2(_09896_),
    .B1(_09897_),
    .X(_09898_));
 sky130_fd_sc_hd__clkbuf_4 _32455_ (.A(_20085_),
    .X(_09899_));
 sky130_fd_sc_hd__nand2_1 _32456_ (.A(_05284_),
    .B(_20081_),
    .Y(_09900_));
 sky130_fd_sc_hd__a21o_1 _32457_ (.A1(_05236_),
    .A2(_09899_),
    .B1(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__buf_6 _32458_ (.A(_09025_),
    .X(_09902_));
 sky130_fd_sc_hd__nand2_1 _32459_ (.A(_05830_),
    .B(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__a21oi_4 _32460_ (.A1(_09898_),
    .A2(_09901_),
    .B1(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__and3_2 _32461_ (.A(_09898_),
    .B(_09901_),
    .C(_09903_),
    .X(_09905_));
 sky130_fd_sc_hd__nor2_8 _32462_ (.A(_09904_),
    .B(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__a21o_1 _32463_ (.A1(_09891_),
    .A2(_09895_),
    .B1(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__nand3_4 _32464_ (.A(_09906_),
    .B(_09891_),
    .C(_09895_),
    .Y(_09908_));
 sky130_fd_sc_hd__o21ai_4 _32465_ (.A1(_09798_),
    .A2(_09784_),
    .B1(_09785_),
    .Y(_09909_));
 sky130_fd_sc_hd__a21o_1 _32466_ (.A1(_09907_),
    .A2(_09908_),
    .B1(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__nand3_4 _32467_ (.A(_09907_),
    .B(_09909_),
    .C(_09908_),
    .Y(_09911_));
 sky130_fd_sc_hd__o21ai_4 _32468_ (.A1(_09788_),
    .A2(_09790_),
    .B1(_09793_),
    .Y(_09912_));
 sky130_fd_sc_hd__a21oi_2 _32469_ (.A1(_09910_),
    .A2(_09911_),
    .B1(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__and3_1 _32470_ (.A(_09907_),
    .B(_09909_),
    .C(_09908_),
    .X(_09914_));
 sky130_fd_sc_hd__nand2_2 _32471_ (.A(_09910_),
    .B(_09912_),
    .Y(_09915_));
 sky130_fd_sc_hd__nor2_2 _32472_ (.A(_09914_),
    .B(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__nand2_1 _32473_ (.A(_09761_),
    .B(_09767_),
    .Y(_09917_));
 sky130_vsdinv _32474_ (.A(_09747_),
    .Y(_09918_));
 sky130_fd_sc_hd__nor2_2 _32475_ (.A(_09750_),
    .B(_09757_),
    .Y(_09919_));
 sky130_fd_sc_hd__nand2_2 _32476_ (.A(_09599_),
    .B(_09600_),
    .Y(_09920_));
 sky130_fd_sc_hd__buf_4 _32477_ (.A(_20114_),
    .X(_09921_));
 sky130_fd_sc_hd__a31o_1 _32478_ (.A1(_09920_),
    .A2(_19910_),
    .A3(_09921_),
    .B1(_09601_),
    .X(_09922_));
 sky130_fd_sc_hd__nand3_4 _32479_ (.A(_06478_),
    .B(_05413_),
    .C(_08057_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_2 _32480_ (.A(_05506_),
    .B(_09476_),
    .Y(_09924_));
 sky130_vsdinv _32481_ (.A(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__buf_4 _32482_ (.A(_08036_),
    .X(_09926_));
 sky130_fd_sc_hd__a22o_1 _32483_ (.A1(_19912_),
    .A2(_08052_),
    .B1(_05608_),
    .B2(_09926_),
    .X(_09927_));
 sky130_fd_sc_hd__o211ai_2 _32484_ (.A1(_08038_),
    .A2(_09923_),
    .B1(_09925_),
    .C1(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__a22oi_4 _32485_ (.A1(_19912_),
    .A2(_08052_),
    .B1(_05608_),
    .B2(_09926_),
    .Y(_09929_));
 sky130_fd_sc_hd__nor2_2 _32486_ (.A(_08037_),
    .B(_09923_),
    .Y(_09930_));
 sky130_fd_sc_hd__o21ai_2 _32487_ (.A1(_09929_),
    .A2(_09930_),
    .B1(_09924_),
    .Y(_09931_));
 sky130_fd_sc_hd__nand3_4 _32488_ (.A(_09922_),
    .B(_09928_),
    .C(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__a21oi_4 _32489_ (.A1(_09603_),
    .A2(_09920_),
    .B1(_09601_),
    .Y(_09933_));
 sky130_fd_sc_hd__o21ai_2 _32490_ (.A1(_09929_),
    .A2(_09930_),
    .B1(_09925_),
    .Y(_09934_));
 sky130_fd_sc_hd__o211ai_4 _32491_ (.A1(_08038_),
    .A2(_09923_),
    .B1(_09924_),
    .C1(_09927_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand3_4 _32492_ (.A(_09933_),
    .B(_09934_),
    .C(_09935_),
    .Y(_09936_));
 sky130_fd_sc_hd__nor2_4 _32493_ (.A(_09740_),
    .B(_09737_),
    .Y(_09937_));
 sky130_vsdinv _32494_ (.A(_09937_),
    .Y(_09938_));
 sky130_fd_sc_hd__a21o_2 _32495_ (.A1(_09932_),
    .A2(_09936_),
    .B1(_09938_),
    .X(_09939_));
 sky130_fd_sc_hd__nand3_4 _32496_ (.A(_09938_),
    .B(_09932_),
    .C(_09936_),
    .Y(_09940_));
 sky130_fd_sc_hd__nand2_1 _32497_ (.A(_09624_),
    .B(_09622_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_4 _32498_ (.A(_09941_),
    .B(_09619_),
    .Y(_09942_));
 sky130_fd_sc_hd__a21oi_4 _32499_ (.A1(_09939_),
    .A2(_09940_),
    .B1(_09942_),
    .Y(_09943_));
 sky130_vsdinv _32500_ (.A(_09932_),
    .Y(_09944_));
 sky130_fd_sc_hd__nand2_1 _32501_ (.A(_09938_),
    .B(_09936_),
    .Y(_09945_));
 sky130_fd_sc_hd__o211a_1 _32502_ (.A1(_09944_),
    .A2(_09945_),
    .B1(_09939_),
    .C1(_09942_),
    .X(_09946_));
 sky130_fd_sc_hd__o22ai_4 _32503_ (.A1(_09918_),
    .A2(_09919_),
    .B1(_09943_),
    .B2(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__a21o_1 _32504_ (.A1(_09939_),
    .A2(_09940_),
    .B1(_09942_),
    .X(_09948_));
 sky130_fd_sc_hd__nand3_4 _32505_ (.A(_09942_),
    .B(_09939_),
    .C(_09940_),
    .Y(_09949_));
 sky130_fd_sc_hd__nand2_2 _32506_ (.A(_09756_),
    .B(_09742_),
    .Y(_09950_));
 sky130_fd_sc_hd__nand3_4 _32507_ (.A(_09948_),
    .B(_09949_),
    .C(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__a22oi_4 _32508_ (.A1(_09766_),
    .A2(_09917_),
    .B1(_09947_),
    .B2(_09951_),
    .Y(_09952_));
 sky130_fd_sc_hd__nor2_1 _32509_ (.A(_09761_),
    .B(_09755_),
    .Y(_09953_));
 sky130_fd_sc_hd__o211a_1 _32510_ (.A1(_09758_),
    .A2(_09953_),
    .B1(_09951_),
    .C1(_09947_),
    .X(_09954_));
 sky130_fd_sc_hd__o22ai_4 _32511_ (.A1(_09913_),
    .A2(_09916_),
    .B1(_09952_),
    .B2(_09954_),
    .Y(_09955_));
 sky130_fd_sc_hd__o21ai_2 _32512_ (.A1(_09761_),
    .A2(_09755_),
    .B1(_09767_),
    .Y(_09956_));
 sky130_fd_sc_hd__a21o_1 _32513_ (.A1(_09947_),
    .A2(_09951_),
    .B1(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__a21oi_1 _32514_ (.A1(_09907_),
    .A2(_09908_),
    .B1(_09909_),
    .Y(_09958_));
 sky130_fd_sc_hd__o21ai_1 _32515_ (.A1(_09958_),
    .A2(_09914_),
    .B1(_09912_),
    .Y(_09959_));
 sky130_fd_sc_hd__nand3b_1 _32516_ (.A_N(_09912_),
    .B(_09910_),
    .C(_09911_),
    .Y(_09960_));
 sky130_fd_sc_hd__nand2_2 _32517_ (.A(_09959_),
    .B(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__nand3_4 _32518_ (.A(_09947_),
    .B(_09956_),
    .C(_09951_),
    .Y(_09962_));
 sky130_fd_sc_hd__nand3_4 _32519_ (.A(_09957_),
    .B(_09961_),
    .C(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__a22oi_4 _32520_ (.A1(_09638_),
    .A2(_09879_),
    .B1(_09955_),
    .B2(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__a21oi_4 _32521_ (.A1(_09636_),
    .A2(_09637_),
    .B1(_09640_),
    .Y(_09965_));
 sky130_fd_sc_hd__o211a_2 _32522_ (.A1(_09634_),
    .A2(_09965_),
    .B1(_09963_),
    .C1(_09955_),
    .X(_09966_));
 sky130_fd_sc_hd__a21bo_1 _32523_ (.A1(_09811_),
    .A2(_09769_),
    .B1_N(_09773_),
    .X(_09967_));
 sky130_fd_sc_hd__o21bai_4 _32524_ (.A1(_09964_),
    .A2(_09966_),
    .B1_N(_09967_),
    .Y(_09968_));
 sky130_vsdinv _32525_ (.A(_09879_),
    .Y(_09969_));
 sky130_fd_sc_hd__o2bb2ai_2 _32526_ (.A1_N(_09963_),
    .A2_N(_09955_),
    .B1(_09632_),
    .B2(_09969_),
    .Y(_09970_));
 sky130_fd_sc_hd__o211ai_4 _32527_ (.A1(_09634_),
    .A2(_09965_),
    .B1(_09963_),
    .C1(_09955_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand3_4 _32528_ (.A(_09970_),
    .B(_09971_),
    .C(_09967_),
    .Y(_09972_));
 sky130_fd_sc_hd__nand2_2 _32529_ (.A(_09968_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__nand3_1 _32530_ (.A(_09729_),
    .B(_09728_),
    .C(_09727_),
    .Y(_09974_));
 sky130_fd_sc_hd__nand2_2 _32531_ (.A(_09974_),
    .B(_09720_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand2_1 _32532_ (.A(_09711_),
    .B(_09713_),
    .Y(_09976_));
 sky130_fd_sc_hd__nand3_4 _32533_ (.A(_19846_),
    .B(_08799_),
    .C(_05243_),
    .Y(_09977_));
 sky130_fd_sc_hd__nor2_8 _32534_ (.A(_05369_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand2_2 _32535_ (.A(\pcpi_mul.rs2[24] ),
    .B(_05289_),
    .Y(_09979_));
 sky130_fd_sc_hd__clkbuf_4 _32536_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09980_));
 sky130_fd_sc_hd__buf_6 _32537_ (.A(_08799_),
    .X(_09981_));
 sky130_fd_sc_hd__a22o_1 _32538_ (.A1(_09980_),
    .A2(_06551_),
    .B1(_09981_),
    .B2(_05549_),
    .X(_09982_));
 sky130_fd_sc_hd__nand3b_4 _32539_ (.A_N(_09978_),
    .B(_09979_),
    .C(_09982_),
    .Y(_09983_));
 sky130_vsdinv _32540_ (.A(_09698_),
    .Y(_09984_));
 sky130_fd_sc_hd__a22oi_4 _32541_ (.A1(_19847_),
    .A2(_06551_),
    .B1(_09981_),
    .B2(_05549_),
    .Y(_09985_));
 sky130_vsdinv _32542_ (.A(_09979_),
    .Y(_09986_));
 sky130_fd_sc_hd__o21ai_2 _32543_ (.A1(_09985_),
    .A2(_09978_),
    .B1(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__nand3_4 _32544_ (.A(_09983_),
    .B(_09984_),
    .C(_09987_),
    .Y(_09988_));
 sky130_fd_sc_hd__nand2_1 _32545_ (.A(_09982_),
    .B(_09986_),
    .Y(_09989_));
 sky130_fd_sc_hd__o21ai_2 _32546_ (.A1(_09985_),
    .A2(_09978_),
    .B1(_09979_),
    .Y(_09990_));
 sky130_fd_sc_hd__o211ai_4 _32547_ (.A1(_09978_),
    .A2(_09989_),
    .B1(_09698_),
    .C1(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__a21oi_1 _32548_ (.A1(_09687_),
    .A2(_09686_),
    .B1(_09681_),
    .Y(_09992_));
 sky130_vsdinv _32549_ (.A(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__a21oi_4 _32550_ (.A1(_09988_),
    .A2(_09991_),
    .B1(_09993_),
    .Y(_09994_));
 sky130_fd_sc_hd__nand2_4 _32551_ (.A(_19843_),
    .B(_05300_),
    .Y(_09995_));
 sky130_fd_sc_hd__buf_4 _32552_ (.A(\pcpi_mul.rs2[29] ),
    .X(_09996_));
 sky130_fd_sc_hd__buf_8 _32553_ (.A(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__clkbuf_8 _32554_ (.A(_19839_),
    .X(_09998_));
 sky130_fd_sc_hd__a22oi_4 _32555_ (.A1(_09997_),
    .A2(_05230_),
    .B1(_09998_),
    .B2(_05418_),
    .Y(_09999_));
 sky130_fd_sc_hd__buf_4 _32556_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10000_));
 sky130_fd_sc_hd__nand2_2 _32557_ (.A(_10000_),
    .B(_05297_),
    .Y(_10001_));
 sky130_fd_sc_hd__nand2_2 _32558_ (.A(_19835_),
    .B(_05214_),
    .Y(_10002_));
 sky130_fd_sc_hd__nor2_4 _32559_ (.A(_10001_),
    .B(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__nor2_4 _32560_ (.A(_09999_),
    .B(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__xnor2_4 _32561_ (.A(_09995_),
    .B(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__nand3_4 _32562_ (.A(_09988_),
    .B(_09991_),
    .C(_09993_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_2 _32563_ (.A(_10005_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__nor2_8 _32564_ (.A(_09994_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__a21o_2 _32565_ (.A1(_09988_),
    .A2(_09991_),
    .B1(_09993_),
    .X(_10009_));
 sky130_fd_sc_hd__a21oi_4 _32566_ (.A1(_10009_),
    .A2(_10006_),
    .B1(_10005_),
    .Y(_10010_));
 sky130_fd_sc_hd__o21ai_4 _32567_ (.A1(_10008_),
    .A2(_10010_),
    .B1(_09703_),
    .Y(_10011_));
 sky130_fd_sc_hd__nand2_2 _32568_ (.A(_10009_),
    .B(_10006_),
    .Y(_10012_));
 sky130_vsdinv _32569_ (.A(_10005_),
    .Y(_10013_));
 sky130_fd_sc_hd__nand2_1 _32570_ (.A(_10012_),
    .B(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__nand3_4 _32571_ (.A(_10009_),
    .B(_10006_),
    .C(_10005_),
    .Y(_10015_));
 sky130_fd_sc_hd__nand3_4 _32572_ (.A(_10014_),
    .B(_09714_),
    .C(_10015_),
    .Y(_10016_));
 sky130_fd_sc_hd__nand2_2 _32573_ (.A(_10011_),
    .B(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__a22oi_4 _32574_ (.A1(_08582_),
    .A2(_05665_),
    .B1(_08775_),
    .B2(_05981_),
    .Y(_10018_));
 sky130_fd_sc_hd__nand3_4 _32575_ (.A(_08315_),
    .B(_19862_),
    .C(_05308_),
    .Y(_10019_));
 sky130_fd_sc_hd__nor2_8 _32576_ (.A(net446),
    .B(_10019_),
    .Y(_10020_));
 sky130_fd_sc_hd__nand2_4 _32577_ (.A(_19865_),
    .B(_06475_),
    .Y(_10021_));
 sky130_vsdinv _32578_ (.A(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__o21ai_2 _32579_ (.A1(_10018_),
    .A2(_10020_),
    .B1(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__a21oi_2 _32580_ (.A1(_09651_),
    .A2(_09648_),
    .B1(_09646_),
    .Y(_10024_));
 sky130_fd_sc_hd__a22o_1 _32581_ (.A1(_08582_),
    .A2(_05665_),
    .B1(_08577_),
    .B2(_05981_),
    .X(_10025_));
 sky130_fd_sc_hd__o211ai_2 _32582_ (.A1(_06256_),
    .A2(_10019_),
    .B1(_10021_),
    .C1(_10025_),
    .Y(_10026_));
 sky130_fd_sc_hd__nand3_4 _32583_ (.A(_10023_),
    .B(_10024_),
    .C(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__nand2_1 _32584_ (.A(_10025_),
    .B(_10022_),
    .Y(_10028_));
 sky130_fd_sc_hd__o22ai_4 _32585_ (.A1(_05580_),
    .A2(_09645_),
    .B1(_09647_),
    .B2(_09644_),
    .Y(_10029_));
 sky130_fd_sc_hd__o21ai_2 _32586_ (.A1(_10018_),
    .A2(_10020_),
    .B1(_10021_),
    .Y(_10030_));
 sky130_fd_sc_hd__o211ai_4 _32587_ (.A1(_10020_),
    .A2(_10028_),
    .B1(_10029_),
    .C1(_10030_),
    .Y(_10031_));
 sky130_fd_sc_hd__nand2_4 _32588_ (.A(_19869_),
    .B(_20148_),
    .Y(_10032_));
 sky130_fd_sc_hd__nand2_4 _32589_ (.A(_07827_),
    .B(_20145_),
    .Y(_10033_));
 sky130_fd_sc_hd__nand2_2 _32590_ (.A(_07356_),
    .B(_06695_),
    .Y(_10034_));
 sky130_fd_sc_hd__a22oi_4 _32591_ (.A1(_08326_),
    .A2(_05827_),
    .B1(_07354_),
    .B2(_07033_),
    .Y(_10035_));
 sky130_fd_sc_hd__nor2_4 _32592_ (.A(_10034_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__o21a_1 _32593_ (.A1(_10032_),
    .A2(_10033_),
    .B1(_10036_),
    .X(_10037_));
 sky130_vsdinv _32594_ (.A(_10034_),
    .Y(_10038_));
 sky130_fd_sc_hd__nor2_8 _32595_ (.A(_10032_),
    .B(_10033_),
    .Y(_10039_));
 sky130_fd_sc_hd__nor2_1 _32596_ (.A(_10035_),
    .B(_10039_),
    .Y(_10040_));
 sky130_fd_sc_hd__nor2_2 _32597_ (.A(_10038_),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__o2bb2ai_4 _32598_ (.A1_N(_10027_),
    .A2_N(_10031_),
    .B1(_10037_),
    .B2(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__nand2_1 _32599_ (.A(_10040_),
    .B(_10034_),
    .Y(_10043_));
 sky130_fd_sc_hd__o21ai_1 _32600_ (.A1(_10035_),
    .A2(_10039_),
    .B1(_10038_),
    .Y(_10044_));
 sky130_fd_sc_hd__nand2_2 _32601_ (.A(_10043_),
    .B(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__nand3_4 _32602_ (.A(_10045_),
    .B(_10031_),
    .C(_10027_),
    .Y(_10046_));
 sky130_vsdinv _32603_ (.A(_09690_),
    .Y(_10047_));
 sky130_fd_sc_hd__a21oi_4 _32604_ (.A1(_10042_),
    .A2(_10046_),
    .B1(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__and3_1 _32605_ (.A(_10042_),
    .B(_10047_),
    .C(_10046_),
    .X(_10049_));
 sky130_fd_sc_hd__nand2_1 _32606_ (.A(_09653_),
    .B(_09670_),
    .Y(_10050_));
 sky130_fd_sc_hd__nand2_4 _32607_ (.A(_10050_),
    .B(_09657_),
    .Y(_10051_));
 sky130_vsdinv _32608_ (.A(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__o21ai_4 _32609_ (.A1(_10048_),
    .A2(_10049_),
    .B1(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__a21o_1 _32610_ (.A1(_10042_),
    .A2(_10046_),
    .B1(_10047_),
    .X(_10054_));
 sky130_fd_sc_hd__nand3_4 _32611_ (.A(_10042_),
    .B(_10047_),
    .C(_10046_),
    .Y(_10055_));
 sky130_fd_sc_hd__nand3_4 _32612_ (.A(_10054_),
    .B(_10055_),
    .C(_10051_),
    .Y(_10056_));
 sky130_fd_sc_hd__nand2_2 _32613_ (.A(_10053_),
    .B(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__nand2_1 _32614_ (.A(_10017_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand2_2 _32615_ (.A(_10015_),
    .B(_09714_),
    .Y(_10059_));
 sky130_fd_sc_hd__o2111ai_4 _32616_ (.A1(_10010_),
    .A2(_10059_),
    .B1(_10056_),
    .C1(_10053_),
    .D1(_10011_),
    .Y(_10060_));
 sky130_fd_sc_hd__nand3_4 _32617_ (.A(_09976_),
    .B(_10058_),
    .C(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__nand3_4 _32618_ (.A(_10017_),
    .B(_10053_),
    .C(_10056_),
    .Y(_10062_));
 sky130_fd_sc_hd__nand3_4 _32619_ (.A(_10057_),
    .B(_10016_),
    .C(_10011_),
    .Y(_10063_));
 sky130_vsdinv _32620_ (.A(_09713_),
    .Y(_10064_));
 sky130_fd_sc_hd__a31oi_4 _32621_ (.A1(_09678_),
    .A2(_09710_),
    .A3(_09715_),
    .B1(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__nand3_4 _32622_ (.A(_10062_),
    .B(_10063_),
    .C(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__buf_6 _32623_ (.A(_07753_),
    .X(_10067_));
 sky130_fd_sc_hd__a22oi_4 _32624_ (.A1(_10067_),
    .A2(_20138_),
    .B1(_07291_),
    .B2(_06442_),
    .Y(_10068_));
 sky130_fd_sc_hd__nand3_4 _32625_ (.A(_19880_),
    .B(_06925_),
    .C(_07028_),
    .Y(_10069_));
 sky130_fd_sc_hd__nor2_4 _32626_ (.A(_06722_),
    .B(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__nand2_2 _32627_ (.A(_07893_),
    .B(_20132_),
    .Y(_10071_));
 sky130_vsdinv _32628_ (.A(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__o21ai_2 _32629_ (.A1(_10068_),
    .A2(_10070_),
    .B1(_10072_),
    .Y(_10073_));
 sky130_fd_sc_hd__a21oi_4 _32630_ (.A1(_09660_),
    .A2(_09662_),
    .B1(_09667_),
    .Y(_10074_));
 sky130_fd_sc_hd__a22o_2 _32631_ (.A1(_07294_),
    .A2(_07502_),
    .B1(_07295_),
    .B2(_06438_),
    .X(_10075_));
 sky130_fd_sc_hd__o211ai_2 _32632_ (.A1(_07510_),
    .A2(_10069_),
    .B1(_10071_),
    .C1(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__nand3_4 _32633_ (.A(_10073_),
    .B(_10074_),
    .C(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__o21ai_2 _32634_ (.A1(_10068_),
    .A2(_10070_),
    .B1(_10071_),
    .Y(_10078_));
 sky130_fd_sc_hd__o21ai_4 _32635_ (.A1(_09661_),
    .A2(_09666_),
    .B1(_09659_),
    .Y(_10079_));
 sky130_fd_sc_hd__o211ai_4 _32636_ (.A1(_07510_),
    .A2(_10069_),
    .B1(_10072_),
    .C1(_10075_),
    .Y(_10080_));
 sky130_fd_sc_hd__nand3_4 _32637_ (.A(_10078_),
    .B(_10079_),
    .C(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__a21o_2 _32638_ (.A1(_09578_),
    .A2(_09579_),
    .B1(_09576_),
    .X(_10082_));
 sky130_fd_sc_hd__a21o_2 _32639_ (.A1(_10077_),
    .A2(_10081_),
    .B1(_10082_),
    .X(_10083_));
 sky130_fd_sc_hd__nand3_4 _32640_ (.A(_10077_),
    .B(_10081_),
    .C(_10082_),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_4 _32641_ (.A(_09595_),
    .B(_09584_),
    .Y(_10085_));
 sky130_fd_sc_hd__a21oi_4 _32642_ (.A1(_10083_),
    .A2(_10084_),
    .B1(_10085_),
    .Y(_10086_));
 sky130_vsdinv _32643_ (.A(_10081_),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_2 _32644_ (.A(_10077_),
    .B(_10082_),
    .Y(_10088_));
 sky130_fd_sc_hd__o211a_2 _32645_ (.A1(_10087_),
    .A2(_10088_),
    .B1(_10083_),
    .C1(_10085_),
    .X(_10089_));
 sky130_fd_sc_hd__nand2_2 _32646_ (.A(_19892_),
    .B(_06713_),
    .Y(_10090_));
 sky130_fd_sc_hd__nand2_2 _32647_ (.A(_06606_),
    .B(_20125_),
    .Y(_10091_));
 sky130_fd_sc_hd__nor2_4 _32648_ (.A(_10090_),
    .B(_10091_),
    .Y(_10092_));
 sky130_vsdinv _32649_ (.A(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__nand2_2 _32650_ (.A(_19898_),
    .B(_06979_),
    .Y(_10094_));
 sky130_vsdinv _32651_ (.A(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__nand2_4 _32652_ (.A(_10090_),
    .B(_10091_),
    .Y(_10096_));
 sky130_fd_sc_hd__nand3_4 _32653_ (.A(_10093_),
    .B(_10095_),
    .C(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__a21o_1 _32654_ (.A1(_09613_),
    .A2(_09614_),
    .B1(_09617_),
    .X(_10098_));
 sky130_fd_sc_hd__a22oi_4 _32655_ (.A1(_19893_),
    .A2(_08151_),
    .B1(_19896_),
    .B2(_20126_),
    .Y(_10099_));
 sky130_fd_sc_hd__o21ai_2 _32656_ (.A1(_10099_),
    .A2(_10092_),
    .B1(_10094_),
    .Y(_10100_));
 sky130_fd_sc_hd__nand3_4 _32657_ (.A(_10097_),
    .B(_10098_),
    .C(_10100_),
    .Y(_10101_));
 sky130_vsdinv _32658_ (.A(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__nand3_2 _32659_ (.A(_10093_),
    .B(_10094_),
    .C(_10096_),
    .Y(_10103_));
 sky130_fd_sc_hd__a21oi_2 _32660_ (.A1(_09613_),
    .A2(_09614_),
    .B1(_09617_),
    .Y(_10104_));
 sky130_fd_sc_hd__o21ai_2 _32661_ (.A1(_10099_),
    .A2(_10092_),
    .B1(_10095_),
    .Y(_10105_));
 sky130_fd_sc_hd__nand3_4 _32662_ (.A(_10103_),
    .B(_10104_),
    .C(_10105_),
    .Y(_10106_));
 sky130_fd_sc_hd__a22oi_4 _32663_ (.A1(_06531_),
    .A2(_07250_),
    .B1(_06196_),
    .B2(_20114_),
    .Y(_10107_));
 sky130_fd_sc_hd__and4_2 _32664_ (.A(_06630_),
    .B(_06534_),
    .C(_07233_),
    .D(_07254_),
    .X(_10108_));
 sky130_fd_sc_hd__nand2_2 _32665_ (.A(_05952_),
    .B(_20110_),
    .Y(_10109_));
 sky130_vsdinv _32666_ (.A(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__o21ai_4 _32667_ (.A1(_10107_),
    .A2(_10108_),
    .B1(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand2_1 _32668_ (.A(_06627_),
    .B(_08042_),
    .Y(_10112_));
 sky130_fd_sc_hd__buf_6 _32669_ (.A(_08433_),
    .X(_10113_));
 sky130_fd_sc_hd__nand3b_4 _32670_ (.A_N(_10112_),
    .B(_06107_),
    .C(_10113_),
    .Y(_10114_));
 sky130_fd_sc_hd__a22o_2 _32671_ (.A1(_06118_),
    .A2(_20118_),
    .B1(_05657_),
    .B2(_07564_),
    .X(_10115_));
 sky130_fd_sc_hd__nand3_4 _32672_ (.A(_10114_),
    .B(_10115_),
    .C(_10109_),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_8 _32673_ (.A(_10111_),
    .B(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__nand2_1 _32674_ (.A(_10106_),
    .B(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__nand2_1 _32675_ (.A(_10101_),
    .B(_10106_),
    .Y(_10119_));
 sky130_vsdinv _32676_ (.A(_10117_),
    .Y(_10120_));
 sky130_fd_sc_hd__nand2_1 _32677_ (.A(_10119_),
    .B(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__o21a_1 _32678_ (.A1(_10102_),
    .A2(_10118_),
    .B1(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__o21ai_1 _32679_ (.A1(_10086_),
    .A2(_10089_),
    .B1(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__a21oi_2 _32680_ (.A1(_09708_),
    .A2(_09676_),
    .B1(_09675_),
    .Y(_10124_));
 sky130_fd_sc_hd__a21o_2 _32681_ (.A1(_10083_),
    .A2(_10084_),
    .B1(_10085_),
    .X(_10125_));
 sky130_fd_sc_hd__nand3_4 _32682_ (.A(_10085_),
    .B(_10083_),
    .C(_10084_),
    .Y(_10126_));
 sky130_fd_sc_hd__nand3_2 _32683_ (.A(_10101_),
    .B(_10106_),
    .C(_10117_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand2_2 _32684_ (.A(_10121_),
    .B(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__nand3_1 _32685_ (.A(_10125_),
    .B(_10126_),
    .C(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand3_2 _32686_ (.A(_10123_),
    .B(_10124_),
    .C(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__clkbuf_4 _32687_ (.A(_10130_),
    .X(_10131_));
 sky130_vsdinv _32688_ (.A(_10127_),
    .Y(_10132_));
 sky130_vsdinv _32689_ (.A(_10121_),
    .Y(_10133_));
 sky130_fd_sc_hd__o22ai_4 _32690_ (.A1(_10132_),
    .A2(_10133_),
    .B1(_10086_),
    .B2(_10089_),
    .Y(_10134_));
 sky130_fd_sc_hd__nand3_4 _32691_ (.A(_10122_),
    .B(_10125_),
    .C(_10126_),
    .Y(_10135_));
 sky130_fd_sc_hd__o21ai_2 _32692_ (.A1(_09677_),
    .A2(_09674_),
    .B1(_09709_),
    .Y(_10136_));
 sky130_fd_sc_hd__nand3_4 _32693_ (.A(_10134_),
    .B(_10135_),
    .C(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2_2 _32694_ (.A(_09630_),
    .B(_09629_),
    .Y(_10138_));
 sky130_fd_sc_hd__clkbuf_4 _32695_ (.A(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__a21oi_4 _32696_ (.A1(_10131_),
    .A2(_10137_),
    .B1(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__and3_1 _32697_ (.A(_10131_),
    .B(_10137_),
    .C(_10139_),
    .X(_10141_));
 sky130_fd_sc_hd__o2bb2ai_2 _32698_ (.A1_N(_10061_),
    .A2_N(_10066_),
    .B1(_10140_),
    .B2(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__and3_2 _32699_ (.A(_10134_),
    .B(_10135_),
    .C(_10136_),
    .X(_10143_));
 sky130_fd_sc_hd__nand2_2 _32700_ (.A(_10130_),
    .B(_10138_),
    .Y(_10144_));
 sky130_fd_sc_hd__nand2_2 _32701_ (.A(_10131_),
    .B(_10137_),
    .Y(_10145_));
 sky130_vsdinv _32702_ (.A(_10139_),
    .Y(_10146_));
 sky130_fd_sc_hd__nand2_4 _32703_ (.A(_10145_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__o2111ai_4 _32704_ (.A1(_10143_),
    .A2(_10144_),
    .B1(_10147_),
    .C1(_10061_),
    .D1(_10066_),
    .Y(_10148_));
 sky130_fd_sc_hd__nand3_4 _32705_ (.A(_09975_),
    .B(_10142_),
    .C(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__nor2_2 _32706_ (.A(_09724_),
    .B(_09726_),
    .Y(_10150_));
 sky130_fd_sc_hd__a31oi_4 _32707_ (.A1(_09729_),
    .A2(_09728_),
    .A3(_09727_),
    .B1(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__o211ai_4 _32708_ (.A1(_10140_),
    .A2(_10141_),
    .B1(_10061_),
    .C1(_10066_),
    .Y(_10152_));
 sky130_fd_sc_hd__a21oi_1 _32709_ (.A1(_10131_),
    .A2(_10137_),
    .B1(_10146_),
    .Y(_10153_));
 sky130_fd_sc_hd__nor2_1 _32710_ (.A(_10139_),
    .B(_10145_),
    .Y(_10154_));
 sky130_fd_sc_hd__o2bb2ai_2 _32711_ (.A1_N(_10061_),
    .A2_N(_10066_),
    .B1(_10153_),
    .B2(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__nand3_4 _32712_ (.A(_10151_),
    .B(_10152_),
    .C(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__nand3_4 _32713_ (.A(_09973_),
    .B(_10149_),
    .C(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__a31oi_4 _32714_ (.A1(_09840_),
    .A2(_09832_),
    .A3(_09818_),
    .B1(_09829_),
    .Y(_10158_));
 sky130_fd_sc_hd__nand2_2 _32715_ (.A(_10156_),
    .B(_10149_),
    .Y(_10159_));
 sky130_fd_sc_hd__nand3_4 _32716_ (.A(_10159_),
    .B(_09972_),
    .C(_09968_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand3_4 _32717_ (.A(_10157_),
    .B(_10158_),
    .C(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_1 _32718_ (.A(_09723_),
    .B(_09730_),
    .Y(_10162_));
 sky130_fd_sc_hd__o22ai_4 _32719_ (.A1(_09838_),
    .A2(_10162_),
    .B1(_09826_),
    .B2(_09833_),
    .Y(_10163_));
 sky130_fd_sc_hd__nand2_1 _32720_ (.A(_09973_),
    .B(_10159_),
    .Y(_10164_));
 sky130_fd_sc_hd__nand2_2 _32721_ (.A(_09970_),
    .B(_09967_),
    .Y(_10165_));
 sky130_fd_sc_hd__o2111ai_4 _32722_ (.A1(_09966_),
    .A2(_10165_),
    .B1(_10149_),
    .C1(_09968_),
    .D1(_10156_),
    .Y(_10166_));
 sky130_fd_sc_hd__nand3_4 _32723_ (.A(_10163_),
    .B(_10164_),
    .C(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand2_1 _32724_ (.A(_10161_),
    .B(_10167_),
    .Y(_10168_));
 sky130_vsdinv _32725_ (.A(_09803_),
    .Y(_10169_));
 sky130_fd_sc_hd__a21oi_4 _32726_ (.A1(_09805_),
    .A2(_09800_),
    .B1(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__a21o_1 _32727_ (.A1(_09818_),
    .A2(_09815_),
    .B1(_10170_),
    .X(_10171_));
 sky130_fd_sc_hd__nand3_2 _32728_ (.A(_09818_),
    .B(_09815_),
    .C(_10170_),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_4 _32729_ (.A(_10171_),
    .B(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nand2_2 _32730_ (.A(_10168_),
    .B(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__a31oi_4 _32731_ (.A1(_10157_),
    .A2(_10158_),
    .A3(_10160_),
    .B1(_10173_),
    .Y(_10175_));
 sky130_fd_sc_hd__nand2_2 _32732_ (.A(_10175_),
    .B(_10167_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand3_4 _32733_ (.A(_09878_),
    .B(_10174_),
    .C(_10176_),
    .Y(_10177_));
 sky130_vsdinv _32734_ (.A(_10173_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand2_1 _32735_ (.A(_10168_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__a21oi_2 _32736_ (.A1(_09819_),
    .A2(_09824_),
    .B1(_09842_),
    .Y(_10180_));
 sky130_fd_sc_hd__a22oi_4 _32737_ (.A1(_10180_),
    .A2(_09834_),
    .B1(_09844_),
    .B2(_09852_),
    .Y(_10181_));
 sky130_fd_sc_hd__nand3_2 _32738_ (.A(_10161_),
    .B(_10167_),
    .C(_10173_),
    .Y(_10182_));
 sky130_fd_sc_hd__nand3_4 _32739_ (.A(_10179_),
    .B(_10181_),
    .C(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__nand2_1 _32740_ (.A(_10177_),
    .B(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__nand2_1 _32741_ (.A(_10184_),
    .B(_09849_),
    .Y(_10185_));
 sky130_vsdinv _32742_ (.A(_09849_),
    .Y(_10186_));
 sky130_fd_sc_hd__nand3_2 _32743_ (.A(_10177_),
    .B(_10183_),
    .C(_10186_),
    .Y(_10187_));
 sky130_fd_sc_hd__a21boi_4 _32744_ (.A1(_09863_),
    .A2(_09865_),
    .B1_N(_09855_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand3_4 _32745_ (.A(_10185_),
    .B(_10187_),
    .C(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__nand2_1 _32746_ (.A(_10184_),
    .B(_10186_),
    .Y(_10190_));
 sky130_fd_sc_hd__nand3_2 _32747_ (.A(_10177_),
    .B(_10183_),
    .C(_09849_),
    .Y(_10191_));
 sky130_fd_sc_hd__nand2_1 _32748_ (.A(_09865_),
    .B(_09863_),
    .Y(_10192_));
 sky130_fd_sc_hd__nand2_1 _32749_ (.A(_10192_),
    .B(_09856_),
    .Y(_10193_));
 sky130_fd_sc_hd__nand3_4 _32750_ (.A(_10190_),
    .B(_10191_),
    .C(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__nand2_2 _32751_ (.A(_10189_),
    .B(_10194_),
    .Y(_10195_));
 sky130_vsdinv _32752_ (.A(_09870_),
    .Y(_10196_));
 sky130_fd_sc_hd__o21ai_4 _32753_ (.A1(_10196_),
    .A2(_09876_),
    .B1(_09867_),
    .Y(_10197_));
 sky130_fd_sc_hd__xor2_4 _32754_ (.A(_10195_),
    .B(_10197_),
    .X(_02648_));
 sky130_fd_sc_hd__a21oi_2 _32755_ (.A1(_09856_),
    .A2(_09865_),
    .B1(_09863_),
    .Y(_10198_));
 sky130_fd_sc_hd__nand2_1 _32756_ (.A(_09869_),
    .B(_09572_),
    .Y(_10199_));
 sky130_fd_sc_hd__o2111ai_4 _32757_ (.A1(_10198_),
    .A2(_10199_),
    .B1(_10189_),
    .C1(_10194_),
    .D1(_09867_),
    .Y(_10200_));
 sky130_vsdinv _32758_ (.A(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand2_1 _32759_ (.A(_09876_),
    .B(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__nand2_1 _32760_ (.A(_10194_),
    .B(_09870_),
    .Y(_10203_));
 sky130_fd_sc_hd__nand2_2 _32761_ (.A(_10203_),
    .B(_10189_),
    .Y(_10204_));
 sky130_fd_sc_hd__a21oi_4 _32762_ (.A1(_10157_),
    .A2(_10160_),
    .B1(_10158_),
    .Y(_10205_));
 sky130_fd_sc_hd__a21oi_4 _32763_ (.A1(_10161_),
    .A2(_10178_),
    .B1(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__nand2_4 _32764_ (.A(_09915_),
    .B(_09911_),
    .Y(_10207_));
 sky130_fd_sc_hd__nand2_4 _32765_ (.A(_10165_),
    .B(_09971_),
    .Y(_10208_));
 sky130_fd_sc_hd__xor2_4 _32766_ (.A(_10207_),
    .B(_10208_),
    .X(_10209_));
 sky130_fd_sc_hd__nand3_1 _32767_ (.A(_09968_),
    .B(_09972_),
    .C(_10156_),
    .Y(_10210_));
 sky130_fd_sc_hd__nand2_2 _32768_ (.A(_10210_),
    .B(_10149_),
    .Y(_10211_));
 sky130_vsdinv _32769_ (.A(_09950_),
    .Y(_10212_));
 sky130_fd_sc_hd__nand2_1 _32770_ (.A(_09949_),
    .B(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__and3_2 _32771_ (.A(_09933_),
    .B(_09934_),
    .C(_09935_),
    .X(_10214_));
 sky130_fd_sc_hd__nor2_2 _32772_ (.A(_09938_),
    .B(_09944_),
    .Y(_10215_));
 sky130_fd_sc_hd__nand3_4 _32773_ (.A(_07660_),
    .B(_06840_),
    .C(_08447_),
    .Y(_10216_));
 sky130_fd_sc_hd__nor2_4 _32774_ (.A(_09047_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__nand2_2 _32775_ (.A(_05506_),
    .B(_20097_),
    .Y(_10218_));
 sky130_fd_sc_hd__a22o_1 _32776_ (.A1(net467),
    .A2(_08884_),
    .B1(_06111_),
    .B2(_08881_),
    .X(_10219_));
 sky130_fd_sc_hd__nand3b_2 _32777_ (.A_N(_10217_),
    .B(_10218_),
    .C(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__a21oi_4 _32778_ (.A1(_10115_),
    .A2(_10110_),
    .B1(_10108_),
    .Y(_10221_));
 sky130_fd_sc_hd__buf_6 _32779_ (.A(_09476_),
    .X(_10222_));
 sky130_fd_sc_hd__a22oi_4 _32780_ (.A1(net467),
    .A2(_08884_),
    .B1(_06111_),
    .B2(_10222_),
    .Y(_10223_));
 sky130_vsdinv _32781_ (.A(_10218_),
    .Y(_10224_));
 sky130_fd_sc_hd__o21ai_2 _32782_ (.A1(_10223_),
    .A2(_10217_),
    .B1(_10224_),
    .Y(_10225_));
 sky130_fd_sc_hd__nand3_4 _32783_ (.A(_10220_),
    .B(_10221_),
    .C(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__o21ai_2 _32784_ (.A1(_10223_),
    .A2(_10217_),
    .B1(_10218_),
    .Y(_10227_));
 sky130_fd_sc_hd__o211ai_2 _32785_ (.A1(_09047_),
    .A2(_10216_),
    .B1(_10224_),
    .C1(_10219_),
    .Y(_10228_));
 sky130_fd_sc_hd__o21ai_2 _32786_ (.A1(_10109_),
    .A2(_10107_),
    .B1(_10114_),
    .Y(_10229_));
 sky130_fd_sc_hd__nand3_4 _32787_ (.A(_10227_),
    .B(_10228_),
    .C(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__nor2_1 _32788_ (.A(_09924_),
    .B(_09929_),
    .Y(_10231_));
 sky130_fd_sc_hd__nor2_1 _32789_ (.A(_09930_),
    .B(_10231_),
    .Y(_10232_));
 sky130_vsdinv _32790_ (.A(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__a21o_2 _32791_ (.A1(_10226_),
    .A2(_10230_),
    .B1(_10233_),
    .X(_10234_));
 sky130_fd_sc_hd__nand3_4 _32792_ (.A(_10233_),
    .B(_10226_),
    .C(_10230_),
    .Y(_10235_));
 sky130_vsdinv _32793_ (.A(_10100_),
    .Y(_10236_));
 sky130_fd_sc_hd__nand2_1 _32794_ (.A(_10097_),
    .B(_10098_),
    .Y(_10237_));
 sky130_fd_sc_hd__o2bb2ai_4 _32795_ (.A1_N(_10106_),
    .A2_N(_10117_),
    .B1(_10236_),
    .B2(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__a21oi_4 _32796_ (.A1(_10234_),
    .A2(_10235_),
    .B1(_10238_),
    .Y(_10239_));
 sky130_vsdinv _32797_ (.A(_10230_),
    .Y(_10240_));
 sky130_fd_sc_hd__nand2_1 _32798_ (.A(_10233_),
    .B(_10226_),
    .Y(_10241_));
 sky130_fd_sc_hd__o211a_2 _32799_ (.A1(_10240_),
    .A2(_10241_),
    .B1(_10234_),
    .C1(_10238_),
    .X(_10242_));
 sky130_fd_sc_hd__o22ai_4 _32800_ (.A1(_10214_),
    .A2(_10215_),
    .B1(_10239_),
    .B2(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__nor2_2 _32801_ (.A(_09937_),
    .B(_10214_),
    .Y(_10244_));
 sky130_fd_sc_hd__nor2_2 _32802_ (.A(_09944_),
    .B(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__nand2_1 _32803_ (.A(_10234_),
    .B(_10235_),
    .Y(_10246_));
 sky130_fd_sc_hd__a21oi_4 _32804_ (.A1(_10106_),
    .A2(_10117_),
    .B1(_10102_),
    .Y(_10247_));
 sky130_fd_sc_hd__nand2_1 _32805_ (.A(_10246_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__nand3_4 _32806_ (.A(_10238_),
    .B(_10234_),
    .C(_10235_),
    .Y(_10249_));
 sky130_fd_sc_hd__nand3b_4 _32807_ (.A_N(_10245_),
    .B(_10248_),
    .C(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__a22oi_4 _32808_ (.A1(_09948_),
    .A2(_10213_),
    .B1(_10243_),
    .B2(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__o2bb2ai_1 _32809_ (.A1_N(_10247_),
    .A2_N(_10246_),
    .B1(_09944_),
    .B2(_10244_),
    .Y(_10252_));
 sky130_fd_sc_hd__o21ai_4 _32810_ (.A1(_10212_),
    .A2(_09943_),
    .B1(_09949_),
    .Y(_10253_));
 sky130_fd_sc_hd__o211a_1 _32811_ (.A1(_10242_),
    .A2(_10252_),
    .B1(_10253_),
    .C1(_10243_),
    .X(_10254_));
 sky130_fd_sc_hd__a21bo_1 _32812_ (.A1(_09906_),
    .A2(_09891_),
    .B1_N(_09895_),
    .X(_10255_));
 sky130_fd_sc_hd__buf_4 _32813_ (.A(\pcpi_mul.rs1[29] ),
    .X(_10256_));
 sky130_fd_sc_hd__nand2_1 _32814_ (.A(_05139_),
    .B(_20081_),
    .Y(_10257_));
 sky130_fd_sc_hd__a21o_1 _32815_ (.A1(_05821_),
    .A2(_10256_),
    .B1(_10257_),
    .X(_10258_));
 sky130_fd_sc_hd__buf_6 _32816_ (.A(\pcpi_mul.rs1[28] ),
    .X(_10259_));
 sky130_fd_sc_hd__nand2_1 _32817_ (.A(_05284_),
    .B(_10256_),
    .Y(_10260_));
 sky130_fd_sc_hd__a21o_1 _32818_ (.A1(_05236_),
    .A2(_10259_),
    .B1(_10260_),
    .X(_10261_));
 sky130_fd_sc_hd__buf_6 _32819_ (.A(_09899_),
    .X(_10262_));
 sky130_fd_sc_hd__nand2_2 _32820_ (.A(_19928_),
    .B(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__a21oi_4 _32821_ (.A1(_10258_),
    .A2(_10261_),
    .B1(_10263_),
    .Y(_10264_));
 sky130_vsdinv _32822_ (.A(_20085_),
    .Y(_10265_));
 sky130_fd_sc_hd__o211a_2 _32823_ (.A1(_05186_),
    .A2(_10265_),
    .B1(_10258_),
    .C1(_10261_),
    .X(_10266_));
 sky130_fd_sc_hd__nor2_8 _32824_ (.A(_10264_),
    .B(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__nand2_2 _32825_ (.A(_05450_),
    .B(_20093_),
    .Y(_10268_));
 sky130_fd_sc_hd__nand2_2 _32826_ (.A(_05312_),
    .B(\pcpi_mul.rs1[26] ),
    .Y(_10269_));
 sky130_fd_sc_hd__nor2_4 _32827_ (.A(_10268_),
    .B(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__and2_1 _32828_ (.A(_10268_),
    .B(_10269_),
    .X(_10271_));
 sky130_fd_sc_hd__nand2_2 _32829_ (.A(_05192_),
    .B(_20072_),
    .Y(_10272_));
 sky130_vsdinv _32830_ (.A(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__o21ai_2 _32831_ (.A1(_10270_),
    .A2(_10271_),
    .B1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__or2_2 _32832_ (.A(_10268_),
    .B(_10269_),
    .X(_10275_));
 sky130_fd_sc_hd__nand2_2 _32833_ (.A(_10268_),
    .B(_10269_),
    .Y(_10276_));
 sky130_fd_sc_hd__nand3_2 _32834_ (.A(_10275_),
    .B(_10272_),
    .C(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__a21oi_4 _32835_ (.A1(_09889_),
    .A2(_09885_),
    .B1(_09887_),
    .Y(_10278_));
 sky130_fd_sc_hd__nand3_4 _32836_ (.A(_10274_),
    .B(_10277_),
    .C(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__o21ai_2 _32837_ (.A1(_10270_),
    .A2(_10271_),
    .B1(_10272_),
    .Y(_10280_));
 sky130_fd_sc_hd__nand3_2 _32838_ (.A(_10275_),
    .B(_10273_),
    .C(_10276_),
    .Y(_10281_));
 sky130_fd_sc_hd__nand3b_4 _32839_ (.A_N(_10278_),
    .B(_10280_),
    .C(_10281_),
    .Y(_10282_));
 sky130_fd_sc_hd__nand3_4 _32840_ (.A(_10267_),
    .B(_10279_),
    .C(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__a21o_1 _32841_ (.A1(_10282_),
    .A2(_10279_),
    .B1(_10267_),
    .X(_10284_));
 sky130_fd_sc_hd__nand3_4 _32842_ (.A(_10255_),
    .B(_10283_),
    .C(_10284_),
    .Y(_10285_));
 sky130_fd_sc_hd__nand2_2 _32843_ (.A(_10284_),
    .B(_10283_),
    .Y(_10286_));
 sky130_fd_sc_hd__a21boi_4 _32844_ (.A1(_09906_),
    .A2(_09891_),
    .B1_N(_09895_),
    .Y(_10287_));
 sky130_fd_sc_hd__o21ba_2 _32845_ (.A1(_09897_),
    .A2(_09900_),
    .B1_N(_09904_),
    .X(_10288_));
 sky130_fd_sc_hd__a21oi_4 _32846_ (.A1(_10286_),
    .A2(_10287_),
    .B1(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__nand2_2 _32847_ (.A(_10286_),
    .B(_10287_),
    .Y(_10290_));
 sky130_fd_sc_hd__a21boi_4 _32848_ (.A1(_10290_),
    .A2(_10285_),
    .B1_N(_10288_),
    .Y(_10291_));
 sky130_fd_sc_hd__a21oi_4 _32849_ (.A1(_10285_),
    .A2(_10289_),
    .B1(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__o21ai_2 _32850_ (.A1(_10251_),
    .A2(_10254_),
    .B1(_10292_),
    .Y(_10293_));
 sky130_fd_sc_hd__a21oi_4 _32851_ (.A1(_10139_),
    .A2(_10131_),
    .B1(_10143_),
    .Y(_10294_));
 sky130_fd_sc_hd__nand2_1 _32852_ (.A(_10290_),
    .B(_10285_),
    .Y(_10295_));
 sky130_fd_sc_hd__nor2_4 _32853_ (.A(_10288_),
    .B(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__nand3_4 _32854_ (.A(_10243_),
    .B(_10253_),
    .C(_10250_),
    .Y(_10297_));
 sky130_fd_sc_hd__a21o_1 _32855_ (.A1(_10243_),
    .A2(_10250_),
    .B1(_10253_),
    .X(_10298_));
 sky130_fd_sc_hd__o211ai_4 _32856_ (.A1(_10291_),
    .A2(_10296_),
    .B1(_10297_),
    .C1(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__nand3_4 _32857_ (.A(_10293_),
    .B(_10294_),
    .C(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__o22ai_2 _32858_ (.A1(_10296_),
    .A2(_10291_),
    .B1(_10251_),
    .B2(_10254_),
    .Y(_10301_));
 sky130_fd_sc_hd__nand3_2 _32859_ (.A(_10298_),
    .B(_10292_),
    .C(_10297_),
    .Y(_10302_));
 sky130_fd_sc_hd__nand2_1 _32860_ (.A(_10144_),
    .B(_10137_),
    .Y(_10303_));
 sky130_fd_sc_hd__nand3_2 _32861_ (.A(_10301_),
    .B(_10302_),
    .C(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__nand2_4 _32862_ (.A(_09963_),
    .B(_09962_),
    .Y(_10305_));
 sky130_fd_sc_hd__a21o_2 _32863_ (.A1(_10300_),
    .A2(_10304_),
    .B1(_10305_),
    .X(_10306_));
 sky130_fd_sc_hd__buf_2 _32864_ (.A(_10304_),
    .X(_10307_));
 sky130_fd_sc_hd__nand3_4 _32865_ (.A(_10300_),
    .B(_10307_),
    .C(_10305_),
    .Y(_10308_));
 sky130_fd_sc_hd__nand2_1 _32866_ (.A(_10306_),
    .B(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand3_4 _32867_ (.A(_10131_),
    .B(_10137_),
    .C(_10139_),
    .Y(_10310_));
 sky130_fd_sc_hd__a21oi_4 _32868_ (.A1(_10062_),
    .A2(_10063_),
    .B1(_10065_),
    .Y(_10311_));
 sky130_fd_sc_hd__a31oi_4 _32869_ (.A1(_10066_),
    .A2(_10147_),
    .A3(_10310_),
    .B1(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__a22oi_4 _32870_ (.A1(_19881_),
    .A2(_06143_),
    .B1(_07090_),
    .B2(_06718_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand3_4 _32871_ (.A(_06927_),
    .B(_07089_),
    .C(_06142_),
    .Y(_10314_));
 sky130_fd_sc_hd__nor2_8 _32872_ (.A(_06440_),
    .B(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__nand2_2 _32873_ (.A(_07893_),
    .B(_06719_),
    .Y(_10316_));
 sky130_fd_sc_hd__o21ai_2 _32874_ (.A1(_10313_),
    .A2(_10315_),
    .B1(_10316_),
    .Y(_10317_));
 sky130_vsdinv _32875_ (.A(_10316_),
    .Y(_10318_));
 sky130_fd_sc_hd__a22o_2 _32876_ (.A1(_19881_),
    .A2(_20135_),
    .B1(_07090_),
    .B2(_06718_),
    .X(_10319_));
 sky130_fd_sc_hd__nand3b_2 _32877_ (.A_N(_10315_),
    .B(_10318_),
    .C(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__o211ai_4 _32878_ (.A1(_10039_),
    .A2(_10036_),
    .B1(_10317_),
    .C1(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__o21ai_2 _32879_ (.A1(_10313_),
    .A2(_10315_),
    .B1(_10318_),
    .Y(_10322_));
 sky130_fd_sc_hd__nand2_1 _32880_ (.A(_10032_),
    .B(_10033_),
    .Y(_10323_));
 sky130_fd_sc_hd__a21oi_4 _32881_ (.A1(_10038_),
    .A2(_10323_),
    .B1(_10039_),
    .Y(_10324_));
 sky130_fd_sc_hd__o211ai_4 _32882_ (.A1(_06452_),
    .A2(_10314_),
    .B1(_10316_),
    .C1(_10319_),
    .Y(_10325_));
 sky130_fd_sc_hd__nand3_4 _32883_ (.A(_10322_),
    .B(_10324_),
    .C(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__a21oi_2 _32884_ (.A1(_10075_),
    .A2(_10072_),
    .B1(_10070_),
    .Y(_10327_));
 sky130_vsdinv _32885_ (.A(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__a21oi_4 _32886_ (.A1(_10321_),
    .A2(_10326_),
    .B1(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__nand3_4 _32887_ (.A(_10321_),
    .B(_10326_),
    .C(_10328_),
    .Y(_10330_));
 sky130_fd_sc_hd__a31o_1 _32888_ (.A1(_10078_),
    .A2(_10079_),
    .A3(_10080_),
    .B1(_10082_),
    .X(_10331_));
 sky130_fd_sc_hd__nand3_2 _32889_ (.A(_10330_),
    .B(_10077_),
    .C(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__nor2_2 _32890_ (.A(_10329_),
    .B(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__a21o_1 _32891_ (.A1(_10321_),
    .A2(_10326_),
    .B1(_10328_),
    .X(_10334_));
 sky130_fd_sc_hd__nand2_4 _32892_ (.A(_10088_),
    .B(_10081_),
    .Y(_10335_));
 sky130_fd_sc_hd__a21oi_2 _32893_ (.A1(_10334_),
    .A2(_10330_),
    .B1(_10335_),
    .Y(_10336_));
 sky130_fd_sc_hd__buf_4 _32894_ (.A(_06531_),
    .X(_10337_));
 sky130_fd_sc_hd__buf_6 _32895_ (.A(_06196_),
    .X(_10338_));
 sky130_fd_sc_hd__a22oi_4 _32896_ (.A1(_10337_),
    .A2(_09921_),
    .B1(_10338_),
    .B2(_20111_),
    .Y(_10339_));
 sky130_fd_sc_hd__buf_6 _32897_ (.A(_09433_),
    .X(_10340_));
 sky130_fd_sc_hd__nand3_4 _32898_ (.A(_06531_),
    .B(_06196_),
    .C(_07561_),
    .Y(_10341_));
 sky130_fd_sc_hd__nor2_4 _32899_ (.A(_10340_),
    .B(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__buf_4 _32900_ (.A(_08057_),
    .X(_10343_));
 sky130_fd_sc_hd__nand2_2 _32901_ (.A(_05953_),
    .B(_10343_),
    .Y(_10344_));
 sky130_vsdinv _32902_ (.A(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__o21ai_2 _32903_ (.A1(_10339_),
    .A2(_10342_),
    .B1(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__buf_4 _32904_ (.A(_06631_),
    .X(_10347_));
 sky130_fd_sc_hd__a22o_1 _32905_ (.A1(_10337_),
    .A2(_09921_),
    .B1(_10347_),
    .B2(_20111_),
    .X(_10348_));
 sky130_fd_sc_hd__nand3b_2 _32906_ (.A_N(_10342_),
    .B(_10348_),
    .C(_10344_),
    .Y(_10349_));
 sky130_fd_sc_hd__clkbuf_4 _32907_ (.A(_07709_),
    .X(_10350_));
 sky130_fd_sc_hd__buf_6 _32908_ (.A(_19896_),
    .X(_10351_));
 sky130_fd_sc_hd__a22oi_2 _32909_ (.A1(_06358_),
    .A2(_10350_),
    .B1(_10351_),
    .B2(_07568_),
    .Y(_10352_));
 sky130_fd_sc_hd__nand2_2 _32910_ (.A(_06357_),
    .B(_08142_),
    .Y(_10353_));
 sky130_fd_sc_hd__nand2_1 _32911_ (.A(_07115_),
    .B(_20123_),
    .Y(_10354_));
 sky130_fd_sc_hd__nor2_1 _32912_ (.A(_10353_),
    .B(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__nand2_2 _32913_ (.A(_19899_),
    .B(_07726_),
    .Y(_10356_));
 sky130_fd_sc_hd__o21bai_2 _32914_ (.A1(_10352_),
    .A2(_10355_),
    .B1_N(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand3b_2 _32915_ (.A_N(_10353_),
    .B(_10351_),
    .C(_20124_),
    .Y(_10358_));
 sky130_fd_sc_hd__nand2_2 _32916_ (.A(_10353_),
    .B(_10354_),
    .Y(_10359_));
 sky130_fd_sc_hd__nand3_4 _32917_ (.A(_10358_),
    .B(_10359_),
    .C(_10356_),
    .Y(_10360_));
 sky130_fd_sc_hd__a21oi_4 _32918_ (.A1(_10095_),
    .A2(_10096_),
    .B1(_10092_),
    .Y(_10361_));
 sky130_fd_sc_hd__a21o_2 _32919_ (.A1(_10357_),
    .A2(_10360_),
    .B1(_10361_),
    .X(_10362_));
 sky130_fd_sc_hd__nand3_4 _32920_ (.A(_10357_),
    .B(_10360_),
    .C(_10361_),
    .Y(_10363_));
 sky130_fd_sc_hd__a22o_1 _32921_ (.A1(_10346_),
    .A2(_10349_),
    .B1(_10362_),
    .B2(_10363_),
    .X(_10364_));
 sky130_fd_sc_hd__nand2_1 _32922_ (.A(_10349_),
    .B(_10346_),
    .Y(_10365_));
 sky130_fd_sc_hd__nand3b_4 _32923_ (.A_N(_10365_),
    .B(_10362_),
    .C(_10363_),
    .Y(_10366_));
 sky130_fd_sc_hd__and2_1 _32924_ (.A(_10364_),
    .B(_10366_),
    .X(_10367_));
 sky130_fd_sc_hd__o21ai_4 _32925_ (.A1(_10333_),
    .A2(_10336_),
    .B1(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__and3_1 _32926_ (.A(_10321_),
    .B(_10326_),
    .C(_10328_),
    .X(_10369_));
 sky130_fd_sc_hd__o21bai_4 _32927_ (.A1(_10329_),
    .A2(_10369_),
    .B1_N(_10335_),
    .Y(_10370_));
 sky130_fd_sc_hd__nand2_4 _32928_ (.A(_10364_),
    .B(_10366_),
    .Y(_10371_));
 sky130_fd_sc_hd__nand3_4 _32929_ (.A(_10334_),
    .B(_10335_),
    .C(_10330_),
    .Y(_10372_));
 sky130_fd_sc_hd__nand3_4 _32930_ (.A(_10370_),
    .B(_10371_),
    .C(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__o21ai_4 _32931_ (.A1(_10052_),
    .A2(_10048_),
    .B1(_10055_),
    .Y(_10374_));
 sky130_fd_sc_hd__a21oi_4 _32932_ (.A1(_10368_),
    .A2(_10373_),
    .B1(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__nand3_4 _32933_ (.A(_10368_),
    .B(_10374_),
    .C(_10373_),
    .Y(_10376_));
 sky130_fd_sc_hd__nand2_2 _32934_ (.A(_10128_),
    .B(_10126_),
    .Y(_10377_));
 sky130_fd_sc_hd__nand2_4 _32935_ (.A(_10377_),
    .B(_10125_),
    .Y(_10378_));
 sky130_fd_sc_hd__nand2_2 _32936_ (.A(_10376_),
    .B(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__nand3_1 _32937_ (.A(_10011_),
    .B(_10053_),
    .C(_10056_),
    .Y(_10380_));
 sky130_fd_sc_hd__nand2_1 _32938_ (.A(_10380_),
    .B(_10016_),
    .Y(_10381_));
 sky130_fd_sc_hd__nor2_2 _32939_ (.A(_09995_),
    .B(_09999_),
    .Y(_10382_));
 sky130_fd_sc_hd__buf_6 _32940_ (.A(_09980_),
    .X(_10383_));
 sky130_fd_sc_hd__buf_6 _32941_ (.A(_19850_),
    .X(_10384_));
 sky130_fd_sc_hd__a22oi_4 _32942_ (.A1(_10383_),
    .A2(_06199_),
    .B1(_10384_),
    .B2(_05481_),
    .Y(_10385_));
 sky130_fd_sc_hd__nor2_4 _32943_ (.A(_09275_),
    .B(_09977_),
    .Y(_10386_));
 sky130_fd_sc_hd__nand2_2 _32944_ (.A(_19853_),
    .B(_05665_),
    .Y(_10387_));
 sky130_fd_sc_hd__o21ai_2 _32945_ (.A1(_10385_),
    .A2(_10386_),
    .B1(_10387_),
    .Y(_10388_));
 sky130_vsdinv _32946_ (.A(_10387_),
    .Y(_10389_));
 sky130_fd_sc_hd__a22o_1 _32947_ (.A1(_10383_),
    .A2(_05244_),
    .B1(_08800_),
    .B2(_05286_),
    .X(_10390_));
 sky130_fd_sc_hd__nand3b_2 _32948_ (.A_N(_10386_),
    .B(_10389_),
    .C(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__o211ai_4 _32949_ (.A1(_10003_),
    .A2(_10382_),
    .B1(_10388_),
    .C1(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__o21ai_4 _32950_ (.A1(_10385_),
    .A2(_10386_),
    .B1(_10389_),
    .Y(_10393_));
 sky130_fd_sc_hd__o21ai_1 _32951_ (.A1(_10001_),
    .A2(_10002_),
    .B1(_09995_),
    .Y(_10394_));
 sky130_fd_sc_hd__nand2_1 _32952_ (.A(_10001_),
    .B(_10002_),
    .Y(_10395_));
 sky130_fd_sc_hd__nand2_2 _32953_ (.A(_10394_),
    .B(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__o211ai_4 _32954_ (.A1(_09275_),
    .A2(_09977_),
    .B1(_10387_),
    .C1(_10390_),
    .Y(_10397_));
 sky130_fd_sc_hd__nand3_4 _32955_ (.A(_10393_),
    .B(_10396_),
    .C(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__nor2_1 _32956_ (.A(_09979_),
    .B(_09985_),
    .Y(_10399_));
 sky130_fd_sc_hd__or2_4 _32957_ (.A(_09978_),
    .B(_10399_),
    .X(_10400_));
 sky130_fd_sc_hd__a21o_2 _32958_ (.A1(_10392_),
    .A2(_10398_),
    .B1(_10400_),
    .X(_10401_));
 sky130_fd_sc_hd__nand3_4 _32959_ (.A(_10400_),
    .B(_10392_),
    .C(_10398_),
    .Y(_10402_));
 sky130_vsdinv _32960_ (.A(_19832_),
    .Y(_10403_));
 sky130_fd_sc_hd__buf_2 _32961_ (.A(_10403_),
    .X(_10404_));
 sky130_fd_sc_hd__buf_8 _32962_ (.A(net441),
    .X(_10405_));
 sky130_fd_sc_hd__nand2_2 _32963_ (.A(_09996_),
    .B(_05131_),
    .Y(_10406_));
 sky130_fd_sc_hd__nand2_2 _32964_ (.A(_10000_),
    .B(_05313_),
    .Y(_10407_));
 sky130_fd_sc_hd__nor2_4 _32965_ (.A(_10406_),
    .B(_10407_),
    .Y(_10408_));
 sky130_fd_sc_hd__nand2_2 _32966_ (.A(_09320_),
    .B(_06614_),
    .Y(_10409_));
 sky130_fd_sc_hd__a21o_1 _32967_ (.A1(_10406_),
    .A2(_10407_),
    .B1(_10409_),
    .X(_10410_));
 sky130_fd_sc_hd__buf_6 _32968_ (.A(_09996_),
    .X(_10411_));
 sky130_fd_sc_hd__buf_8 _32969_ (.A(_19839_),
    .X(_10412_));
 sky130_fd_sc_hd__a22oi_4 _32970_ (.A1(_10411_),
    .A2(_07901_),
    .B1(_10412_),
    .B2(_06197_),
    .Y(_10413_));
 sky130_fd_sc_hd__o21ai_2 _32971_ (.A1(_10413_),
    .A2(_10408_),
    .B1(_10409_),
    .Y(_10414_));
 sky130_fd_sc_hd__o21ai_1 _32972_ (.A1(_10408_),
    .A2(_10410_),
    .B1(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__o21ai_2 _32973_ (.A1(_10405_),
    .A2(_04840_),
    .B1(_10415_),
    .Y(_10416_));
 sky130_fd_sc_hd__nor2_2 _32974_ (.A(_10404_),
    .B(_04839_),
    .Y(_10417_));
 sky130_fd_sc_hd__o211ai_4 _32975_ (.A1(_10408_),
    .A2(_10410_),
    .B1(_10417_),
    .C1(_10414_),
    .Y(_10418_));
 sky130_fd_sc_hd__nand2_4 _32976_ (.A(_10416_),
    .B(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__a21boi_4 _32977_ (.A1(_10401_),
    .A2(_10402_),
    .B1_N(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__a21oi_2 _32978_ (.A1(_10392_),
    .A2(_10398_),
    .B1(_10400_),
    .Y(_10421_));
 sky130_fd_sc_hd__nor3b_4 _32979_ (.A(_10419_),
    .B(_10421_),
    .C_N(_10402_),
    .Y(_10422_));
 sky130_fd_sc_hd__o22ai_4 _32980_ (.A1(_10013_),
    .A2(_10012_),
    .B1(_10420_),
    .B2(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__nand2_1 _32981_ (.A(_10401_),
    .B(_10402_),
    .Y(_10424_));
 sky130_fd_sc_hd__nand2_2 _32982_ (.A(_10424_),
    .B(_10419_),
    .Y(_10425_));
 sky130_fd_sc_hd__nand3b_4 _32983_ (.A_N(_10419_),
    .B(_10402_),
    .C(_10401_),
    .Y(_10426_));
 sky130_fd_sc_hd__nand3_4 _32984_ (.A(_10425_),
    .B(_10008_),
    .C(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__nand2_1 _32985_ (.A(_10423_),
    .B(_10427_),
    .Y(_10428_));
 sky130_vsdinv _32986_ (.A(_10027_),
    .Y(_10429_));
 sky130_fd_sc_hd__and3_1 _32987_ (.A(_10031_),
    .B(_10044_),
    .C(_10043_),
    .X(_10430_));
 sky130_fd_sc_hd__nand3_4 _32988_ (.A(_08589_),
    .B(_08575_),
    .C(_05799_),
    .Y(_10431_));
 sky130_fd_sc_hd__nor2_8 _32989_ (.A(_08243_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__buf_6 _32990_ (.A(_08773_),
    .X(_10433_));
 sky130_fd_sc_hd__a22o_2 _32991_ (.A1(_10433_),
    .A2(_05573_),
    .B1(_07965_),
    .B2(_20152_),
    .X(_10434_));
 sky130_fd_sc_hd__buf_8 _32992_ (.A(\pcpi_mul.rs2[21] ),
    .X(_10435_));
 sky130_fd_sc_hd__nand2_4 _32993_ (.A(_10435_),
    .B(_06480_),
    .Y(_10436_));
 sky130_vsdinv _32994_ (.A(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_1 _32995_ (.A(_10434_),
    .B(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__o22ai_4 _32996_ (.A1(_06256_),
    .A2(_10019_),
    .B1(_10021_),
    .B2(_10018_),
    .Y(_10439_));
 sky130_fd_sc_hd__buf_8 _32997_ (.A(_08773_),
    .X(_10440_));
 sky130_fd_sc_hd__a22oi_4 _32998_ (.A1(_10440_),
    .A2(_05693_),
    .B1(_19863_),
    .B2(_05991_),
    .Y(_10441_));
 sky130_fd_sc_hd__o21ai_2 _32999_ (.A1(_10441_),
    .A2(_10432_),
    .B1(_10436_),
    .Y(_10442_));
 sky130_fd_sc_hd__o211ai_4 _33000_ (.A1(_10432_),
    .A2(_10438_),
    .B1(_10439_),
    .C1(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__o21ai_2 _33001_ (.A1(_10441_),
    .A2(_10432_),
    .B1(_10437_),
    .Y(_10444_));
 sky130_fd_sc_hd__a21oi_2 _33002_ (.A1(_10025_),
    .A2(_10022_),
    .B1(_10020_),
    .Y(_10445_));
 sky130_fd_sc_hd__buf_6 _33003_ (.A(_08242_),
    .X(_10446_));
 sky130_fd_sc_hd__o211ai_4 _33004_ (.A1(_10446_),
    .A2(_10431_),
    .B1(_10436_),
    .C1(_10434_),
    .Y(_10447_));
 sky130_fd_sc_hd__nand3_4 _33005_ (.A(_10444_),
    .B(_10445_),
    .C(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__nand2_4 _33006_ (.A(_08326_),
    .B(_05826_),
    .Y(_10449_));
 sky130_fd_sc_hd__nand2_4 _33007_ (.A(_19873_),
    .B(_07024_),
    .Y(_10450_));
 sky130_fd_sc_hd__nor2_8 _33008_ (.A(_10449_),
    .B(_10450_),
    .Y(_10451_));
 sky130_fd_sc_hd__and2_1 _33009_ (.A(_10449_),
    .B(_10450_),
    .X(_10452_));
 sky130_fd_sc_hd__nand2_2 _33010_ (.A(_19877_),
    .B(_05986_),
    .Y(_10453_));
 sky130_vsdinv _33011_ (.A(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__o21ai_2 _33012_ (.A1(_10451_),
    .A2(_10452_),
    .B1(_10454_),
    .Y(_10455_));
 sky130_fd_sc_hd__nand2_2 _33013_ (.A(_10449_),
    .B(_10450_),
    .Y(_10456_));
 sky130_fd_sc_hd__nand3b_4 _33014_ (.A_N(_10451_),
    .B(_10456_),
    .C(_10453_),
    .Y(_10457_));
 sky130_fd_sc_hd__nand2_4 _33015_ (.A(_10455_),
    .B(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__a21o_1 _33016_ (.A1(_10443_),
    .A2(_10448_),
    .B1(_10458_),
    .X(_10459_));
 sky130_fd_sc_hd__nand3_4 _33017_ (.A(_10458_),
    .B(_10443_),
    .C(_10448_),
    .Y(_10460_));
 sky130_fd_sc_hd__a21oi_1 _33018_ (.A1(_09983_),
    .A2(_09987_),
    .B1(_09984_),
    .Y(_10461_));
 sky130_fd_sc_hd__a21o_1 _33019_ (.A1(_09988_),
    .A2(_09993_),
    .B1(_10461_),
    .X(_10462_));
 sky130_fd_sc_hd__a21oi_4 _33020_ (.A1(_10459_),
    .A2(_10460_),
    .B1(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__a21oi_4 _33021_ (.A1(_10443_),
    .A2(_10448_),
    .B1(_10458_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_1 _33022_ (.A(_09991_),
    .B(_09992_),
    .Y(_10465_));
 sky130_fd_sc_hd__nand2_2 _33023_ (.A(_10465_),
    .B(_09988_),
    .Y(_10466_));
 sky130_fd_sc_hd__nor3_1 _33024_ (.A(_10454_),
    .B(_10451_),
    .C(_10452_),
    .Y(_10467_));
 sky130_fd_sc_hd__o21a_1 _33025_ (.A1(_10451_),
    .A2(_10452_),
    .B1(_10454_),
    .X(_10468_));
 sky130_fd_sc_hd__o211a_2 _33026_ (.A1(_10467_),
    .A2(_10468_),
    .B1(_10448_),
    .C1(_10443_),
    .X(_10469_));
 sky130_fd_sc_hd__nor3_4 _33027_ (.A(_10464_),
    .B(_10466_),
    .C(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__o22ai_4 _33028_ (.A1(_10429_),
    .A2(_10430_),
    .B1(_10463_),
    .B2(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__o21ai_4 _33029_ (.A1(_10464_),
    .A2(_10469_),
    .B1(_10466_),
    .Y(_10472_));
 sky130_fd_sc_hd__nand3_4 _33030_ (.A(_10462_),
    .B(_10460_),
    .C(_10459_),
    .Y(_10473_));
 sky130_fd_sc_hd__nand2_1 _33031_ (.A(_10045_),
    .B(_10027_),
    .Y(_10474_));
 sky130_fd_sc_hd__nand2_4 _33032_ (.A(_10474_),
    .B(_10031_),
    .Y(_10475_));
 sky130_fd_sc_hd__nand3_4 _33033_ (.A(_10472_),
    .B(_10473_),
    .C(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__nand2_1 _33034_ (.A(_10471_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__nand2_2 _33035_ (.A(_10428_),
    .B(_10477_),
    .Y(_10478_));
 sky130_fd_sc_hd__nand2_2 _33036_ (.A(_10008_),
    .B(_10426_),
    .Y(_10479_));
 sky130_fd_sc_hd__o2111ai_4 _33037_ (.A1(_10420_),
    .A2(_10479_),
    .B1(_10476_),
    .C1(_10471_),
    .D1(_10423_),
    .Y(_10480_));
 sky130_fd_sc_hd__nand3_4 _33038_ (.A(_10381_),
    .B(_10478_),
    .C(_10480_),
    .Y(_10481_));
 sky130_fd_sc_hd__nand3_2 _33039_ (.A(_10428_),
    .B(_10476_),
    .C(_10471_),
    .Y(_10482_));
 sky130_fd_sc_hd__nor2_2 _33040_ (.A(_10010_),
    .B(_10059_),
    .Y(_10483_));
 sky130_fd_sc_hd__a31oi_4 _33041_ (.A1(_10011_),
    .A2(_10053_),
    .A3(_10056_),
    .B1(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__nand3_2 _33042_ (.A(_10477_),
    .B(_10427_),
    .C(_10423_),
    .Y(_10485_));
 sky130_fd_sc_hd__nand3_4 _33043_ (.A(_10482_),
    .B(_10484_),
    .C(_10485_),
    .Y(_10486_));
 sky130_fd_sc_hd__nand2_1 _33044_ (.A(_10052_),
    .B(_10055_),
    .Y(_10487_));
 sky130_fd_sc_hd__nand2_2 _33045_ (.A(_10487_),
    .B(_10054_),
    .Y(_10488_));
 sky130_fd_sc_hd__a21oi_4 _33046_ (.A1(_10370_),
    .A2(_10372_),
    .B1(_10371_),
    .Y(_10489_));
 sky130_fd_sc_hd__o211a_2 _33047_ (.A1(_10329_),
    .A2(_10332_),
    .B1(_10371_),
    .C1(_10370_),
    .X(_10490_));
 sky130_fd_sc_hd__nor3_4 _33048_ (.A(_10488_),
    .B(_10489_),
    .C(_10490_),
    .Y(_10491_));
 sky130_vsdinv _33049_ (.A(_10378_),
    .Y(_10492_));
 sky130_fd_sc_hd__o21ai_2 _33050_ (.A1(_10375_),
    .A2(_10491_),
    .B1(_10492_),
    .Y(_10493_));
 sky130_fd_sc_hd__o2111ai_4 _33051_ (.A1(_10375_),
    .A2(_10379_),
    .B1(_10481_),
    .C1(_10486_),
    .D1(_10493_),
    .Y(_10494_));
 sky130_vsdinv _33052_ (.A(_10487_),
    .Y(_10495_));
 sky130_fd_sc_hd__o22ai_4 _33053_ (.A1(_10048_),
    .A2(_10495_),
    .B1(_10489_),
    .B2(_10490_),
    .Y(_10496_));
 sky130_fd_sc_hd__a21oi_1 _33054_ (.A1(_10496_),
    .A2(_10376_),
    .B1(_10378_),
    .Y(_10497_));
 sky130_fd_sc_hd__nor2_1 _33055_ (.A(_10375_),
    .B(_10379_),
    .Y(_10498_));
 sky130_fd_sc_hd__o2bb2ai_2 _33056_ (.A1_N(_10481_),
    .A2_N(_10486_),
    .B1(_10497_),
    .B2(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__nand3_4 _33057_ (.A(_10312_),
    .B(_10494_),
    .C(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__nand3_1 _33058_ (.A(_10066_),
    .B(_10147_),
    .C(_10310_),
    .Y(_10501_));
 sky130_fd_sc_hd__nand2_2 _33059_ (.A(_10501_),
    .B(_10061_),
    .Y(_10502_));
 sky130_fd_sc_hd__a21oi_1 _33060_ (.A1(_10496_),
    .A2(_10376_),
    .B1(_10492_),
    .Y(_10503_));
 sky130_fd_sc_hd__nor2_1 _33061_ (.A(_10128_),
    .B(_10086_),
    .Y(_10504_));
 sky130_fd_sc_hd__o211a_1 _33062_ (.A1(_10089_),
    .A2(_10504_),
    .B1(_10376_),
    .C1(_10496_),
    .X(_10505_));
 sky130_fd_sc_hd__o2bb2ai_2 _33063_ (.A1_N(_10481_),
    .A2_N(_10486_),
    .B1(_10503_),
    .B2(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__nand2_2 _33064_ (.A(_10496_),
    .B(_10492_),
    .Y(_10507_));
 sky130_vsdinv _33065_ (.A(_10377_),
    .Y(_10508_));
 sky130_fd_sc_hd__o22ai_4 _33066_ (.A1(_10086_),
    .A2(_10508_),
    .B1(_10375_),
    .B2(_10491_),
    .Y(_10509_));
 sky130_fd_sc_hd__o2111ai_4 _33067_ (.A1(_10491_),
    .A2(_10507_),
    .B1(_10481_),
    .C1(_10486_),
    .D1(_10509_),
    .Y(_10510_));
 sky130_fd_sc_hd__nand3_4 _33068_ (.A(_10502_),
    .B(_10506_),
    .C(_10510_),
    .Y(_10511_));
 sky130_fd_sc_hd__nand2_1 _33069_ (.A(_10500_),
    .B(_10511_),
    .Y(_10512_));
 sky130_fd_sc_hd__nand2_2 _33070_ (.A(_10309_),
    .B(_10512_),
    .Y(_10513_));
 sky130_fd_sc_hd__nand2_2 _33071_ (.A(_10300_),
    .B(_10305_),
    .Y(_10514_));
 sky130_vsdinv _33072_ (.A(_10307_),
    .Y(_10515_));
 sky130_fd_sc_hd__o2111ai_4 _33073_ (.A1(_10514_),
    .A2(_10515_),
    .B1(_10511_),
    .C1(_10500_),
    .D1(_10306_),
    .Y(_10516_));
 sky130_fd_sc_hd__nand3_4 _33074_ (.A(_10211_),
    .B(_10513_),
    .C(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__a21oi_2 _33075_ (.A1(_10152_),
    .A2(_10155_),
    .B1(_10151_),
    .Y(_10518_));
 sky130_fd_sc_hd__a31oi_4 _33076_ (.A1(_09968_),
    .A2(_10156_),
    .A3(_09972_),
    .B1(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__nand3_2 _33077_ (.A(_10512_),
    .B(_10308_),
    .C(_10306_),
    .Y(_10520_));
 sky130_fd_sc_hd__a21oi_2 _33078_ (.A1(_10300_),
    .A2(_10307_),
    .B1(_10305_),
    .Y(_10521_));
 sky130_fd_sc_hd__and2_1 _33079_ (.A(_09957_),
    .B(_09961_),
    .X(_10522_));
 sky130_fd_sc_hd__o211a_1 _33080_ (.A1(_09954_),
    .A2(_10522_),
    .B1(_10307_),
    .C1(_10300_),
    .X(_10523_));
 sky130_fd_sc_hd__o211ai_4 _33081_ (.A1(_10521_),
    .A2(_10523_),
    .B1(_10511_),
    .C1(_10500_),
    .Y(_10524_));
 sky130_fd_sc_hd__nand3_4 _33082_ (.A(_10519_),
    .B(_10520_),
    .C(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__nand3b_2 _33083_ (.A_N(_10209_),
    .B(_10517_),
    .C(_10525_),
    .Y(_10526_));
 sky130_vsdinv _33084_ (.A(_10208_),
    .Y(_10527_));
 sky130_fd_sc_hd__nor2_1 _33085_ (.A(_10207_),
    .B(_10527_),
    .Y(_10528_));
 sky130_vsdinv _33086_ (.A(_10207_),
    .Y(_10529_));
 sky130_fd_sc_hd__nor2_1 _33087_ (.A(_10529_),
    .B(_10208_),
    .Y(_10530_));
 sky130_fd_sc_hd__o2bb2ai_2 _33088_ (.A1_N(_10525_),
    .A2_N(_10517_),
    .B1(_10528_),
    .B2(_10530_),
    .Y(_10531_));
 sky130_fd_sc_hd__nand3_4 _33089_ (.A(_10206_),
    .B(_10526_),
    .C(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__nand3_4 _33090_ (.A(_10209_),
    .B(_10517_),
    .C(_10525_),
    .Y(_10533_));
 sky130_fd_sc_hd__nor2_4 _33091_ (.A(_10529_),
    .B(_10527_),
    .Y(_10534_));
 sky130_fd_sc_hd__nor2_1 _33092_ (.A(_10207_),
    .B(_10208_),
    .Y(_10535_));
 sky130_fd_sc_hd__o2bb2ai_2 _33093_ (.A1_N(_10525_),
    .A2_N(_10517_),
    .B1(_10534_),
    .B2(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__o211ai_4 _33094_ (.A1(_10205_),
    .A2(_10175_),
    .B1(_10533_),
    .C1(_10536_),
    .Y(_10537_));
 sky130_vsdinv _33095_ (.A(_10171_),
    .Y(_10538_));
 sky130_fd_sc_hd__a21oi_1 _33096_ (.A1(_10532_),
    .A2(_10537_),
    .B1(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__and3_1 _33097_ (.A(_10532_),
    .B(_10537_),
    .C(_10538_),
    .X(_10540_));
 sky130_vsdinv _33098_ (.A(_10176_),
    .Y(_10541_));
 sky130_fd_sc_hd__nand2_1 _33099_ (.A(_09878_),
    .B(_10174_),
    .Y(_10542_));
 sky130_fd_sc_hd__o2bb2ai_2 _33100_ (.A1_N(_09849_),
    .A2_N(_10183_),
    .B1(_10541_),
    .B2(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__o21bai_2 _33101_ (.A1(_10539_),
    .A2(_10540_),
    .B1_N(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__nand2_1 _33102_ (.A(_10532_),
    .B(_10538_),
    .Y(_10545_));
 sky130_vsdinv _33103_ (.A(_10537_),
    .Y(_10546_));
 sky130_fd_sc_hd__a21o_1 _33104_ (.A1(_10532_),
    .A2(_10537_),
    .B1(_10538_),
    .X(_10547_));
 sky130_fd_sc_hd__o211ai_4 _33105_ (.A1(_10545_),
    .A2(_10546_),
    .B1(_10543_),
    .C1(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__nand2_1 _33106_ (.A(_10544_),
    .B(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__a21oi_1 _33107_ (.A1(_10202_),
    .A2(_10204_),
    .B1(_10549_),
    .Y(_10550_));
 sky130_fd_sc_hd__and3_1 _33108_ (.A(_10202_),
    .B(_10549_),
    .C(_10204_),
    .X(_10551_));
 sky130_fd_sc_hd__nor2_1 _33109_ (.A(_10550_),
    .B(_10551_),
    .Y(_02649_));
 sky130_fd_sc_hd__buf_6 _33110_ (.A(_09980_),
    .X(_10552_));
 sky130_fd_sc_hd__buf_6 _33111_ (.A(_19850_),
    .X(_10553_));
 sky130_fd_sc_hd__a22oi_4 _33112_ (.A1(_10552_),
    .A2(_06348_),
    .B1(_10553_),
    .B2(_05675_),
    .Y(_10554_));
 sky130_fd_sc_hd__nand3_4 _33113_ (.A(_19847_),
    .B(_09981_),
    .C(_20162_),
    .Y(_10555_));
 sky130_fd_sc_hd__nor2_4 _33114_ (.A(_05580_),
    .B(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__nand2_2 _33115_ (.A(_08802_),
    .B(_05981_),
    .Y(_10557_));
 sky130_fd_sc_hd__o21ai_2 _33116_ (.A1(_10554_),
    .A2(_10556_),
    .B1(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__nand3b_1 _33117_ (.A_N(_10406_),
    .B(_19841_),
    .C(_05144_),
    .Y(_10559_));
 sky130_fd_sc_hd__o21ai_2 _33118_ (.A1(_10409_),
    .A2(_10413_),
    .B1(_10559_),
    .Y(_10560_));
 sky130_vsdinv _33119_ (.A(_10557_),
    .Y(_10561_));
 sky130_fd_sc_hd__a22o_4 _33120_ (.A1(_10383_),
    .A2(_05867_),
    .B1(_10384_),
    .B2(_05474_),
    .X(_10562_));
 sky130_fd_sc_hd__o211ai_4 _33121_ (.A1(_05296_),
    .A2(_10555_),
    .B1(_10561_),
    .C1(_10562_),
    .Y(_10563_));
 sky130_fd_sc_hd__and3_2 _33122_ (.A(_10558_),
    .B(_10560_),
    .C(_10563_),
    .X(_10564_));
 sky130_fd_sc_hd__o21ai_2 _33123_ (.A1(_10554_),
    .A2(_10556_),
    .B1(_10561_),
    .Y(_10565_));
 sky130_fd_sc_hd__o21ai_1 _33124_ (.A1(_10406_),
    .A2(_10407_),
    .B1(_10409_),
    .Y(_10566_));
 sky130_fd_sc_hd__nand2_1 _33125_ (.A(_10406_),
    .B(_10407_),
    .Y(_10567_));
 sky130_fd_sc_hd__nand2_1 _33126_ (.A(_10566_),
    .B(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__o211ai_2 _33127_ (.A1(_05296_),
    .A2(_10555_),
    .B1(_10557_),
    .C1(_10562_),
    .Y(_10569_));
 sky130_fd_sc_hd__nand3_4 _33128_ (.A(_10565_),
    .B(_10568_),
    .C(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__a21o_2 _33129_ (.A1(_10390_),
    .A2(_10389_),
    .B1(_10386_),
    .X(_10571_));
 sky130_fd_sc_hd__nand2_4 _33130_ (.A(_10570_),
    .B(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__clkbuf_8 _33131_ (.A(_19832_),
    .X(_10573_));
 sky130_fd_sc_hd__a22oi_4 _33132_ (.A1(_19829_),
    .A2(_05230_),
    .B1(_10573_),
    .B2(_20174_),
    .Y(_10574_));
 sky130_fd_sc_hd__buf_6 _33133_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10575_));
 sky130_fd_sc_hd__nand2_2 _33134_ (.A(_10575_),
    .B(_04838_),
    .Y(_10576_));
 sky130_fd_sc_hd__clkbuf_8 _33135_ (.A(\pcpi_mul.rs2[30] ),
    .X(_10577_));
 sky130_fd_sc_hd__nand2_2 _33136_ (.A(_10577_),
    .B(_05417_),
    .Y(_10578_));
 sky130_fd_sc_hd__nor2_8 _33137_ (.A(_10576_),
    .B(_10578_),
    .Y(_10579_));
 sky130_fd_sc_hd__nand2_4 _33138_ (.A(\pcpi_mul.rs2[29] ),
    .B(_20170_),
    .Y(_10580_));
 sky130_fd_sc_hd__nand3b_4 _33139_ (.A_N(_10580_),
    .B(_09998_),
    .C(_05177_),
    .Y(_10581_));
 sky130_fd_sc_hd__nand2_4 _33140_ (.A(_10000_),
    .B(_06551_),
    .Y(_10582_));
 sky130_fd_sc_hd__nand2_2 _33141_ (.A(_10580_),
    .B(_10582_),
    .Y(_10583_));
 sky130_fd_sc_hd__nand2_4 _33142_ (.A(_09696_),
    .B(_05549_),
    .Y(_10584_));
 sky130_fd_sc_hd__nand3_4 _33143_ (.A(_10581_),
    .B(_10583_),
    .C(_10584_),
    .Y(_10585_));
 sky130_fd_sc_hd__a22oi_4 _33144_ (.A1(_10411_),
    .A2(_20171_),
    .B1(_10412_),
    .B2(_06614_),
    .Y(_10586_));
 sky130_fd_sc_hd__nor2_4 _33145_ (.A(_10580_),
    .B(_10582_),
    .Y(_10587_));
 sky130_vsdinv _33146_ (.A(_10584_),
    .Y(_10588_));
 sky130_fd_sc_hd__o21ai_2 _33147_ (.A1(_10586_),
    .A2(_10587_),
    .B1(_10588_),
    .Y(_10589_));
 sky130_fd_sc_hd__o211ai_4 _33148_ (.A1(_10574_),
    .A2(_10579_),
    .B1(_10585_),
    .C1(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__o21ai_2 _33149_ (.A1(_10586_),
    .A2(_10587_),
    .B1(_10584_),
    .Y(_10591_));
 sky130_fd_sc_hd__a21oi_4 _33150_ (.A1(_10580_),
    .A2(_10582_),
    .B1(_10584_),
    .Y(_10592_));
 sky130_fd_sc_hd__nand2_1 _33151_ (.A(_10592_),
    .B(_10581_),
    .Y(_10593_));
 sky130_fd_sc_hd__nor2_2 _33152_ (.A(_10574_),
    .B(_10579_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand3_4 _33153_ (.A(_10591_),
    .B(_10593_),
    .C(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__nand3b_4 _33154_ (.A_N(_10418_),
    .B(_10590_),
    .C(_10595_),
    .Y(_10596_));
 sky130_fd_sc_hd__nand2_1 _33155_ (.A(_10590_),
    .B(_10595_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_4 _33156_ (.A(_10597_),
    .B(_10418_),
    .Y(_10598_));
 sky130_fd_sc_hd__nand3_4 _33157_ (.A(_10558_),
    .B(_10560_),
    .C(_10563_),
    .Y(_10599_));
 sky130_fd_sc_hd__a21o_1 _33158_ (.A1(_10570_),
    .A2(_10599_),
    .B1(_10571_),
    .X(_10600_));
 sky130_fd_sc_hd__o2111ai_4 _33159_ (.A1(_10564_),
    .A2(_10572_),
    .B1(_10596_),
    .C1(_10598_),
    .D1(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__a21oi_2 _33160_ (.A1(_10599_),
    .A2(_10570_),
    .B1(_10571_),
    .Y(_10602_));
 sky130_fd_sc_hd__nor2_2 _33161_ (.A(_10564_),
    .B(_10572_),
    .Y(_10603_));
 sky130_fd_sc_hd__o2bb2ai_4 _33162_ (.A1_N(_10596_),
    .A2_N(_10598_),
    .B1(_10602_),
    .B2(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__o2bb2ai_2 _33163_ (.A1_N(_10601_),
    .A2_N(_10604_),
    .B1(_10419_),
    .B2(_10424_),
    .Y(_10605_));
 sky130_fd_sc_hd__nand3_4 _33164_ (.A(_10422_),
    .B(_10604_),
    .C(_10601_),
    .Y(_10606_));
 sky130_fd_sc_hd__nand2_1 _33165_ (.A(_10605_),
    .B(_10606_),
    .Y(_10607_));
 sky130_vsdinv _33166_ (.A(_10448_),
    .Y(_10608_));
 sky130_fd_sc_hd__and3_1 _33167_ (.A(_10443_),
    .B(_10455_),
    .C(_10457_),
    .X(_10609_));
 sky130_fd_sc_hd__buf_4 _33168_ (.A(_08773_),
    .X(_10610_));
 sky130_fd_sc_hd__buf_4 _33169_ (.A(_05555_),
    .X(_10611_));
 sky130_fd_sc_hd__a22oi_4 _33170_ (.A1(_10610_),
    .A2(_06476_),
    .B1(_08592_),
    .B2(_10611_),
    .Y(_10612_));
 sky130_fd_sc_hd__nand3_4 _33171_ (.A(_08773_),
    .B(_08591_),
    .C(_06480_),
    .Y(_10613_));
 sky130_fd_sc_hd__nor2_4 _33172_ (.A(_08243_),
    .B(_10613_),
    .Y(_10614_));
 sky130_fd_sc_hd__nand2_4 _33173_ (.A(_10435_),
    .B(_06841_),
    .Y(_10615_));
 sky130_vsdinv _33174_ (.A(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__o21ai_2 _33175_ (.A1(_10612_),
    .A2(_10614_),
    .B1(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__a21oi_2 _33176_ (.A1(_10434_),
    .A2(_10437_),
    .B1(_10432_),
    .Y(_10618_));
 sky130_fd_sc_hd__buf_4 _33177_ (.A(_10613_),
    .X(_10619_));
 sky130_fd_sc_hd__buf_6 _33178_ (.A(_19862_),
    .X(_10620_));
 sky130_fd_sc_hd__a22o_2 _33179_ (.A1(_10610_),
    .A2(_20152_),
    .B1(_10620_),
    .B2(_10611_),
    .X(_10621_));
 sky130_fd_sc_hd__o211ai_4 _33180_ (.A1(_10446_),
    .A2(_10619_),
    .B1(_10615_),
    .C1(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__nand3_4 _33181_ (.A(_10617_),
    .B(_10618_),
    .C(_10622_),
    .Y(_10623_));
 sky130_fd_sc_hd__o21ai_2 _33182_ (.A1(_10612_),
    .A2(_10614_),
    .B1(_10615_),
    .Y(_10624_));
 sky130_fd_sc_hd__o211ai_4 _33183_ (.A1(_10446_),
    .A2(_10619_),
    .B1(_10616_),
    .C1(_10621_),
    .Y(_10625_));
 sky130_fd_sc_hd__o22ai_4 _33184_ (.A1(_10446_),
    .A2(_10431_),
    .B1(_10436_),
    .B2(_10441_),
    .Y(_10626_));
 sky130_fd_sc_hd__nand3_4 _33185_ (.A(_10624_),
    .B(_10625_),
    .C(_10626_),
    .Y(_10627_));
 sky130_fd_sc_hd__buf_4 _33186_ (.A(_19869_),
    .X(_10628_));
 sky130_fd_sc_hd__a22oi_4 _33187_ (.A1(_10628_),
    .A2(_05999_),
    .B1(_07973_),
    .B2(_05986_),
    .Y(_10629_));
 sky130_fd_sc_hd__nand2_2 _33188_ (.A(_08779_),
    .B(_06695_),
    .Y(_10630_));
 sky130_fd_sc_hd__nand2_2 _33189_ (.A(_08598_),
    .B(_06696_),
    .Y(_10631_));
 sky130_fd_sc_hd__nor2_4 _33190_ (.A(_10630_),
    .B(_10631_),
    .Y(_10632_));
 sky130_fd_sc_hd__nor2_1 _33191_ (.A(_10629_),
    .B(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__nand2_2 _33192_ (.A(_19877_),
    .B(_06442_),
    .Y(_10634_));
 sky130_fd_sc_hd__nand2_1 _33193_ (.A(_10633_),
    .B(_10634_),
    .Y(_10635_));
 sky130_vsdinv _33194_ (.A(_10634_),
    .Y(_10636_));
 sky130_fd_sc_hd__o21ai_2 _33195_ (.A1(_10629_),
    .A2(_10632_),
    .B1(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__nand2_4 _33196_ (.A(_10635_),
    .B(_10637_),
    .Y(_10638_));
 sky130_fd_sc_hd__a21o_2 _33197_ (.A1(_10623_),
    .A2(_10627_),
    .B1(_10638_),
    .X(_10639_));
 sky130_fd_sc_hd__nand3_4 _33198_ (.A(_10638_),
    .B(_10627_),
    .C(_10623_),
    .Y(_10640_));
 sky130_fd_sc_hd__a21oi_4 _33199_ (.A1(_10393_),
    .A2(_10397_),
    .B1(_10396_),
    .Y(_10641_));
 sky130_fd_sc_hd__a21o_2 _33200_ (.A1(_10400_),
    .A2(_10398_),
    .B1(_10641_),
    .X(_10642_));
 sky130_fd_sc_hd__a21oi_4 _33201_ (.A1(_10639_),
    .A2(_10640_),
    .B1(_10642_),
    .Y(_10643_));
 sky130_fd_sc_hd__o21a_1 _33202_ (.A1(_09978_),
    .A2(_10399_),
    .B1(_10398_),
    .X(_10644_));
 sky130_fd_sc_hd__o211a_2 _33203_ (.A1(_10641_),
    .A2(_10644_),
    .B1(_10640_),
    .C1(_10639_),
    .X(_10645_));
 sky130_fd_sc_hd__o22ai_4 _33204_ (.A1(_10608_),
    .A2(_10609_),
    .B1(_10643_),
    .B2(_10645_),
    .Y(_10646_));
 sky130_fd_sc_hd__a21oi_2 _33205_ (.A1(_10623_),
    .A2(_10627_),
    .B1(_10638_),
    .Y(_10647_));
 sky130_fd_sc_hd__nor3_2 _33206_ (.A(_10636_),
    .B(_10629_),
    .C(_10632_),
    .Y(_10648_));
 sky130_fd_sc_hd__nor2_1 _33207_ (.A(_10634_),
    .B(_10633_),
    .Y(_10649_));
 sky130_fd_sc_hd__o211a_1 _33208_ (.A1(_10648_),
    .A2(_10649_),
    .B1(_10627_),
    .C1(_10623_),
    .X(_10650_));
 sky130_fd_sc_hd__nor2_2 _33209_ (.A(_10641_),
    .B(_10644_),
    .Y(_10651_));
 sky130_fd_sc_hd__o21ai_4 _33210_ (.A1(_10647_),
    .A2(_10650_),
    .B1(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__nand3_4 _33211_ (.A(_10642_),
    .B(_10639_),
    .C(_10640_),
    .Y(_10653_));
 sky130_fd_sc_hd__nand2_1 _33212_ (.A(_10458_),
    .B(_10448_),
    .Y(_10654_));
 sky130_fd_sc_hd__nand2_2 _33213_ (.A(_10654_),
    .B(_10443_),
    .Y(_10655_));
 sky130_fd_sc_hd__nand3_4 _33214_ (.A(_10652_),
    .B(_10653_),
    .C(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__nand2_1 _33215_ (.A(_10646_),
    .B(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand2_4 _33216_ (.A(_10607_),
    .B(_10657_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand2_1 _33217_ (.A(_10652_),
    .B(_10655_),
    .Y(_10659_));
 sky130_fd_sc_hd__o2111ai_4 _33218_ (.A1(_10645_),
    .A2(_10659_),
    .B1(_10606_),
    .C1(_10646_),
    .D1(_10605_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand2_1 _33219_ (.A(_10658_),
    .B(_10660_),
    .Y(_10661_));
 sky130_fd_sc_hd__nand3_2 _33220_ (.A(_10423_),
    .B(_10471_),
    .C(_10476_),
    .Y(_10662_));
 sky130_fd_sc_hd__o21a_1 _33221_ (.A1(_10420_),
    .A2(_10479_),
    .B1(_10662_),
    .X(_10663_));
 sky130_fd_sc_hd__nand2_2 _33222_ (.A(_10661_),
    .B(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__nand2_2 _33223_ (.A(_10662_),
    .B(_10427_),
    .Y(_10665_));
 sky130_fd_sc_hd__nand3_4 _33224_ (.A(_10665_),
    .B(_10658_),
    .C(_10660_),
    .Y(_10666_));
 sky130_fd_sc_hd__nand2_1 _33225_ (.A(_10664_),
    .B(_10666_),
    .Y(_10667_));
 sky130_fd_sc_hd__nand3_4 _33226_ (.A(_10067_),
    .B(_07295_),
    .C(_08002_),
    .Y(_10668_));
 sky130_fd_sc_hd__a22o_2 _33227_ (.A1(_07289_),
    .A2(_20133_),
    .B1(_07291_),
    .B2(_08151_),
    .X(_10669_));
 sky130_fd_sc_hd__o21ai_1 _33228_ (.A1(_06452_),
    .A2(_10668_),
    .B1(_10669_),
    .Y(_10670_));
 sky130_fd_sc_hd__nand2_2 _33229_ (.A(_19890_),
    .B(_20126_),
    .Y(_10671_));
 sky130_vsdinv _33230_ (.A(_10671_),
    .Y(_10672_));
 sky130_fd_sc_hd__nand2_2 _33231_ (.A(_10670_),
    .B(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__a21oi_4 _33232_ (.A1(_10454_),
    .A2(_10456_),
    .B1(_10451_),
    .Y(_10674_));
 sky130_fd_sc_hd__o211ai_4 _33233_ (.A1(_06452_),
    .A2(_10668_),
    .B1(_10671_),
    .C1(_10669_),
    .Y(_10675_));
 sky130_fd_sc_hd__nand3_4 _33234_ (.A(_10673_),
    .B(_10674_),
    .C(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__nand2_1 _33235_ (.A(_10670_),
    .B(_10671_),
    .Y(_10677_));
 sky130_fd_sc_hd__nor2_4 _33236_ (.A(_06440_),
    .B(_10668_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand3b_4 _33237_ (.A_N(_10678_),
    .B(_10672_),
    .C(_10669_),
    .Y(_10679_));
 sky130_fd_sc_hd__nand3b_4 _33238_ (.A_N(_10674_),
    .B(_10677_),
    .C(_10679_),
    .Y(_10680_));
 sky130_fd_sc_hd__nor2_2 _33239_ (.A(_10318_),
    .B(_10315_),
    .Y(_10681_));
 sky130_fd_sc_hd__o2bb2ai_4 _33240_ (.A1_N(_10676_),
    .A2_N(_10680_),
    .B1(_10313_),
    .B2(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__a21oi_4 _33241_ (.A1(_10319_),
    .A2(_10318_),
    .B1(_10315_),
    .Y(_10683_));
 sky130_fd_sc_hd__a31oi_4 _33242_ (.A1(_10673_),
    .A2(_10674_),
    .A3(_10675_),
    .B1(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__nand2_4 _33243_ (.A(_10684_),
    .B(_10680_),
    .Y(_10685_));
 sky130_fd_sc_hd__nand2_4 _33244_ (.A(_10330_),
    .B(_10321_),
    .Y(_10686_));
 sky130_fd_sc_hd__a21oi_4 _33245_ (.A1(_10682_),
    .A2(_10685_),
    .B1(_10686_),
    .Y(_10687_));
 sky130_fd_sc_hd__a31oi_1 _33246_ (.A1(_10322_),
    .A2(_10324_),
    .A3(_10325_),
    .B1(_10327_),
    .Y(_10688_));
 sky130_vsdinv _33247_ (.A(_10321_),
    .Y(_10689_));
 sky130_fd_sc_hd__o211a_2 _33248_ (.A1(_10688_),
    .A2(_10689_),
    .B1(_10685_),
    .C1(_10682_),
    .X(_10690_));
 sky130_fd_sc_hd__buf_6 _33249_ (.A(_07718_),
    .X(_10691_));
 sky130_fd_sc_hd__buf_4 _33250_ (.A(_07922_),
    .X(_10692_));
 sky130_fd_sc_hd__buf_6 _33251_ (.A(_06207_),
    .X(_10693_));
 sky130_fd_sc_hd__buf_4 _33252_ (.A(_07251_),
    .X(_10694_));
 sky130_fd_sc_hd__nand3_4 _33253_ (.A(_10692_),
    .B(_10693_),
    .C(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand2_1 _33254_ (.A(_06544_),
    .B(_06976_),
    .Y(_10696_));
 sky130_fd_sc_hd__nand2_1 _33255_ (.A(_19896_),
    .B(_20118_),
    .Y(_10697_));
 sky130_fd_sc_hd__nand2_2 _33256_ (.A(_10696_),
    .B(_10697_),
    .Y(_10698_));
 sky130_fd_sc_hd__o21ai_1 _33257_ (.A1(_10691_),
    .A2(_10695_),
    .B1(_10698_),
    .Y(_10699_));
 sky130_fd_sc_hd__buf_4 _33258_ (.A(_07785_),
    .X(_10700_));
 sky130_fd_sc_hd__nand2_2 _33259_ (.A(_10700_),
    .B(_07561_),
    .Y(_10701_));
 sky130_vsdinv _33260_ (.A(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__nand2_2 _33261_ (.A(_10699_),
    .B(_10702_),
    .Y(_10703_));
 sky130_fd_sc_hd__buf_6 _33262_ (.A(_07718_),
    .X(_10704_));
 sky130_fd_sc_hd__o211ai_4 _33263_ (.A1(_10704_),
    .A2(_10695_),
    .B1(_10701_),
    .C1(_10698_),
    .Y(_10705_));
 sky130_fd_sc_hd__o21ai_1 _33264_ (.A1(_10353_),
    .A2(_10354_),
    .B1(_10356_),
    .Y(_10706_));
 sky130_fd_sc_hd__nand2_2 _33265_ (.A(_10706_),
    .B(_10359_),
    .Y(_10707_));
 sky130_fd_sc_hd__a21o_1 _33266_ (.A1(_10703_),
    .A2(_10705_),
    .B1(_10707_),
    .X(_10708_));
 sky130_vsdinv _33267_ (.A(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__nand3_4 _33268_ (.A(_10703_),
    .B(_10707_),
    .C(_10705_),
    .Y(_10710_));
 sky130_fd_sc_hd__buf_4 _33269_ (.A(_20110_),
    .X(_10711_));
 sky130_fd_sc_hd__a22oi_4 _33270_ (.A1(_06119_),
    .A2(_10711_),
    .B1(_10347_),
    .B2(_10343_),
    .Y(_10712_));
 sky130_fd_sc_hd__nand2_2 _33271_ (.A(_06118_),
    .B(_08053_),
    .Y(_10713_));
 sky130_fd_sc_hd__nand2_1 _33272_ (.A(_06107_),
    .B(_08453_),
    .Y(_10714_));
 sky130_fd_sc_hd__nor2_1 _33273_ (.A(_10713_),
    .B(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__buf_4 _33274_ (.A(_08447_),
    .X(_10716_));
 sky130_fd_sc_hd__nand2_2 _33275_ (.A(_05953_),
    .B(_10716_),
    .Y(_10717_));
 sky130_fd_sc_hd__o21bai_1 _33276_ (.A1(_10712_),
    .A2(_10715_),
    .B1_N(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__nand3b_2 _33277_ (.A_N(_10713_),
    .B(_10338_),
    .C(_20108_),
    .Y(_10719_));
 sky130_fd_sc_hd__nand2_1 _33278_ (.A(_10713_),
    .B(_10714_),
    .Y(_10720_));
 sky130_fd_sc_hd__nand3_1 _33279_ (.A(_10719_),
    .B(_10717_),
    .C(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__nand2_2 _33280_ (.A(_10718_),
    .B(_10721_),
    .Y(_10722_));
 sky130_fd_sc_hd__nand2_2 _33281_ (.A(_10710_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__a21o_1 _33282_ (.A1(_10708_),
    .A2(_10710_),
    .B1(_10722_),
    .X(_10724_));
 sky130_fd_sc_hd__o21ai_4 _33283_ (.A1(_10709_),
    .A2(_10723_),
    .B1(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__o21ai_2 _33284_ (.A1(_10687_),
    .A2(_10690_),
    .B1(_10725_),
    .Y(_10726_));
 sky130_vsdinv _33285_ (.A(_10475_),
    .Y(_10727_));
 sky130_fd_sc_hd__o21ai_4 _33286_ (.A1(_10727_),
    .A2(_10463_),
    .B1(_10473_),
    .Y(_10728_));
 sky130_fd_sc_hd__o21a_1 _33287_ (.A1(_10709_),
    .A2(_10723_),
    .B1(_10724_),
    .X(_10729_));
 sky130_fd_sc_hd__a21o_1 _33288_ (.A1(_10682_),
    .A2(_10685_),
    .B1(_10686_),
    .X(_10730_));
 sky130_fd_sc_hd__nand3_4 _33289_ (.A(_10686_),
    .B(_10682_),
    .C(_10685_),
    .Y(_10731_));
 sky130_fd_sc_hd__nand3_4 _33290_ (.A(_10729_),
    .B(_10730_),
    .C(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__nand3_4 _33291_ (.A(_10726_),
    .B(_10728_),
    .C(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__nand2_1 _33292_ (.A(_10708_),
    .B(_10710_),
    .Y(_10734_));
 sky130_fd_sc_hd__nor2_2 _33293_ (.A(_10722_),
    .B(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__and2_1 _33294_ (.A(_10734_),
    .B(_10722_),
    .X(_10736_));
 sky130_fd_sc_hd__o22ai_4 _33295_ (.A1(_10735_),
    .A2(_10736_),
    .B1(_10687_),
    .B2(_10690_),
    .Y(_10737_));
 sky130_fd_sc_hd__a21oi_4 _33296_ (.A1(_10472_),
    .A2(_10475_),
    .B1(_10470_),
    .Y(_10738_));
 sky130_fd_sc_hd__nand3_2 _33297_ (.A(_10730_),
    .B(_10731_),
    .C(_10725_),
    .Y(_10739_));
 sky130_fd_sc_hd__nand3_4 _33298_ (.A(_10737_),
    .B(_10738_),
    .C(_10739_),
    .Y(_10740_));
 sky130_fd_sc_hd__a21o_2 _33299_ (.A1(_10370_),
    .A2(_10371_),
    .B1(_10333_),
    .X(_10741_));
 sky130_fd_sc_hd__a21o_2 _33300_ (.A1(_10733_),
    .A2(_10740_),
    .B1(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__nand3_4 _33301_ (.A(_10733_),
    .B(_10740_),
    .C(_10741_),
    .Y(_10743_));
 sky130_fd_sc_hd__nand2_2 _33302_ (.A(_10742_),
    .B(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__nand2_2 _33303_ (.A(_10667_),
    .B(_10744_),
    .Y(_10745_));
 sky130_fd_sc_hd__o211ai_4 _33304_ (.A1(_10491_),
    .A2(_10507_),
    .B1(_10486_),
    .C1(_10509_),
    .Y(_10746_));
 sky130_fd_sc_hd__nand2_4 _33305_ (.A(_10746_),
    .B(_10481_),
    .Y(_10747_));
 sky130_vsdinv _33306_ (.A(_10733_),
    .Y(_10748_));
 sky130_fd_sc_hd__nand2_1 _33307_ (.A(_10740_),
    .B(_10741_),
    .Y(_10749_));
 sky130_fd_sc_hd__o2111ai_4 _33308_ (.A1(_10748_),
    .A2(_10749_),
    .B1(_10742_),
    .C1(_10666_),
    .D1(_10664_),
    .Y(_10750_));
 sky130_fd_sc_hd__nand3_4 _33309_ (.A(_10745_),
    .B(_10747_),
    .C(_10750_),
    .Y(_10751_));
 sky130_fd_sc_hd__a22oi_4 _33310_ (.A1(_10742_),
    .A2(_10743_),
    .B1(_10664_),
    .B2(_10666_),
    .Y(_10752_));
 sky130_fd_sc_hd__a21oi_4 _33311_ (.A1(_10658_),
    .A2(_10660_),
    .B1(_10665_),
    .Y(_10753_));
 sky130_fd_sc_hd__nand3_2 _33312_ (.A(_10666_),
    .B(_10742_),
    .C(_10743_),
    .Y(_10754_));
 sky130_fd_sc_hd__nor2_2 _33313_ (.A(_10753_),
    .B(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__nand2_1 _33314_ (.A(_10478_),
    .B(_10480_),
    .Y(_10756_));
 sky130_fd_sc_hd__o21a_1 _33315_ (.A1(_10484_),
    .A2(_10756_),
    .B1(_10746_),
    .X(_10757_));
 sky130_fd_sc_hd__o21ai_4 _33316_ (.A1(_10752_),
    .A2(_10755_),
    .B1(_10757_),
    .Y(_10758_));
 sky130_fd_sc_hd__a21bo_1 _33317_ (.A1(_10279_),
    .A2(_10267_),
    .B1_N(_10282_),
    .X(_10759_));
 sky130_fd_sc_hd__buf_4 _33318_ (.A(_20072_),
    .X(_10760_));
 sky130_fd_sc_hd__buf_4 _33319_ (.A(_20077_),
    .X(_10761_));
 sky130_fd_sc_hd__and4_2 _33320_ (.A(_05140_),
    .B(_05142_),
    .C(_10760_),
    .D(_10761_),
    .X(_10762_));
 sky130_fd_sc_hd__buf_8 _33321_ (.A(_09775_),
    .X(_10763_));
 sky130_fd_sc_hd__nor2_4 _33322_ (.A(_05154_),
    .B(_10763_),
    .Y(_10764_));
 sky130_vsdinv _33323_ (.A(_10764_),
    .Y(_10765_));
 sky130_vsdinv _33324_ (.A(\pcpi_mul.rs1[30] ),
    .Y(_10766_));
 sky130_fd_sc_hd__clkbuf_8 _33325_ (.A(_10766_),
    .X(_10767_));
 sky130_fd_sc_hd__buf_6 _33326_ (.A(_20077_),
    .X(_10768_));
 sky130_fd_sc_hd__nand2_2 _33327_ (.A(_19932_),
    .B(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__o21ai_4 _33328_ (.A1(_05151_),
    .A2(_10767_),
    .B1(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__nand3b_4 _33329_ (.A_N(_10762_),
    .B(_10765_),
    .C(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__buf_6 _33330_ (.A(_10766_),
    .X(_10772_));
 sky130_fd_sc_hd__o21a_1 _33331_ (.A1(_05151_),
    .A2(_10772_),
    .B1(_10769_),
    .X(_10773_));
 sky130_fd_sc_hd__o21ai_4 _33332_ (.A1(_10762_),
    .A2(_10773_),
    .B1(_10764_),
    .Y(_10774_));
 sky130_fd_sc_hd__nand2_8 _33333_ (.A(_10771_),
    .B(_10774_),
    .Y(_10775_));
 sky130_vsdinv _33334_ (.A(_10775_),
    .Y(_10776_));
 sky130_fd_sc_hd__buf_4 _33335_ (.A(\pcpi_mul.rs1[31] ),
    .X(_10777_));
 sky130_fd_sc_hd__buf_6 _33336_ (.A(_10777_),
    .X(_10778_));
 sky130_fd_sc_hd__buf_6 _33337_ (.A(_10778_),
    .X(_10779_));
 sky130_vsdinv _33338_ (.A(\pcpi_mul.rs1[26] ),
    .Y(_10780_));
 sky130_fd_sc_hd__buf_6 _33339_ (.A(_10780_),
    .X(_10781_));
 sky130_fd_sc_hd__nand3_2 _33340_ (.A(_19921_),
    .B(_05805_),
    .C(_09787_),
    .Y(_10782_));
 sky130_fd_sc_hd__nand2_1 _33341_ (.A(_05816_),
    .B(_20090_),
    .Y(_10783_));
 sky130_fd_sc_hd__nand2_2 _33342_ (.A(_05674_),
    .B(_09474_),
    .Y(_10784_));
 sky130_fd_sc_hd__nand2_2 _33343_ (.A(_10783_),
    .B(_10784_),
    .Y(_10785_));
 sky130_fd_sc_hd__o21ai_2 _33344_ (.A1(_10781_),
    .A2(_10782_),
    .B1(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__a21o_1 _33345_ (.A1(_19939_),
    .A2(_10779_),
    .B1(_10786_),
    .X(_10787_));
 sky130_fd_sc_hd__nand2_2 _33346_ (.A(_19938_),
    .B(_10778_),
    .Y(_10788_));
 sky130_vsdinv _33347_ (.A(_10788_),
    .Y(_10789_));
 sky130_fd_sc_hd__nand2_1 _33348_ (.A(_10786_),
    .B(_10789_),
    .Y(_10790_));
 sky130_fd_sc_hd__a21oi_4 _33349_ (.A1(_10273_),
    .A2(_10276_),
    .B1(_10270_),
    .Y(_10791_));
 sky130_fd_sc_hd__nand3_4 _33350_ (.A(_10787_),
    .B(_10790_),
    .C(_10791_),
    .Y(_10792_));
 sky130_fd_sc_hd__nor2_1 _33351_ (.A(_10783_),
    .B(_10784_),
    .Y(_10793_));
 sky130_fd_sc_hd__nand3b_2 _33352_ (.A_N(_10793_),
    .B(_10785_),
    .C(_10789_),
    .Y(_10794_));
 sky130_fd_sc_hd__nand2_1 _33353_ (.A(_10786_),
    .B(_10788_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand3b_4 _33354_ (.A_N(_10791_),
    .B(_10794_),
    .C(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand2_1 _33355_ (.A(_10792_),
    .B(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__nand2_1 _33356_ (.A(_10776_),
    .B(_10797_),
    .Y(_10798_));
 sky130_fd_sc_hd__nand3_2 _33357_ (.A(_10792_),
    .B(_10775_),
    .C(_10796_),
    .Y(_10799_));
 sky130_fd_sc_hd__nand3_4 _33358_ (.A(_10759_),
    .B(_10798_),
    .C(_10799_),
    .Y(_10800_));
 sky130_fd_sc_hd__nand3_2 _33359_ (.A(_10776_),
    .B(_10796_),
    .C(_10792_),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_1 _33360_ (.A(_10797_),
    .B(_10775_),
    .Y(_10802_));
 sky130_fd_sc_hd__a21boi_2 _33361_ (.A1(_10267_),
    .A2(_10279_),
    .B1_N(_10282_),
    .Y(_10803_));
 sky130_fd_sc_hd__nand3_4 _33362_ (.A(_10801_),
    .B(_10802_),
    .C(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__nor2_1 _33363_ (.A(_10257_),
    .B(_10260_),
    .Y(_10805_));
 sky130_fd_sc_hd__or2_2 _33364_ (.A(_10805_),
    .B(_10264_),
    .X(_10806_));
 sky130_fd_sc_hd__a21oi_4 _33365_ (.A1(_10800_),
    .A2(_10804_),
    .B1(_10806_),
    .Y(_10807_));
 sky130_fd_sc_hd__and3_2 _33366_ (.A(_10800_),
    .B(_10804_),
    .C(_10806_),
    .X(_10808_));
 sky130_fd_sc_hd__clkbuf_4 _33367_ (.A(_05502_),
    .X(_10809_));
 sky130_fd_sc_hd__a22oi_4 _33368_ (.A1(_10809_),
    .A2(_09044_),
    .B1(_19916_),
    .B2(_20098_),
    .Y(_10810_));
 sky130_fd_sc_hd__buf_4 _33369_ (.A(_09476_),
    .X(_10811_));
 sky130_fd_sc_hd__nand3_4 _33370_ (.A(_06096_),
    .B(_05414_),
    .C(_10811_),
    .Y(_10812_));
 sky130_fd_sc_hd__nor2_4 _33371_ (.A(_08888_),
    .B(_10812_),
    .Y(_10813_));
 sky130_fd_sc_hd__buf_4 _33372_ (.A(_20093_),
    .X(_10814_));
 sky130_fd_sc_hd__nand2_2 _33373_ (.A(_19918_),
    .B(_10814_),
    .Y(_10815_));
 sky130_vsdinv _33374_ (.A(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__o21ai_2 _33375_ (.A1(_10810_),
    .A2(_10813_),
    .B1(_10816_),
    .Y(_10817_));
 sky130_fd_sc_hd__a21oi_4 _33376_ (.A1(_10348_),
    .A2(_10345_),
    .B1(_10342_),
    .Y(_10818_));
 sky130_fd_sc_hd__a22o_2 _33377_ (.A1(_19913_),
    .A2(_20102_),
    .B1(_19916_),
    .B2(_20098_),
    .X(_10819_));
 sky130_fd_sc_hd__o211ai_4 _33378_ (.A1(_09880_),
    .A2(_10812_),
    .B1(_10815_),
    .C1(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__nand3_4 _33379_ (.A(_10817_),
    .B(_10818_),
    .C(_10820_),
    .Y(_10821_));
 sky130_fd_sc_hd__o21ai_2 _33380_ (.A1(_10810_),
    .A2(_10813_),
    .B1(_10815_),
    .Y(_10822_));
 sky130_fd_sc_hd__o211ai_4 _33381_ (.A1(_09880_),
    .A2(_10812_),
    .B1(_10816_),
    .C1(_10819_),
    .Y(_10823_));
 sky130_fd_sc_hd__buf_4 _33382_ (.A(_10340_),
    .X(_10824_));
 sky130_fd_sc_hd__o22ai_4 _33383_ (.A1(_10824_),
    .A2(_10341_),
    .B1(_10344_),
    .B2(_10339_),
    .Y(_10825_));
 sky130_fd_sc_hd__nand3_4 _33384_ (.A(_10822_),
    .B(_10823_),
    .C(_10825_),
    .Y(_10826_));
 sky130_fd_sc_hd__nor2_4 _33385_ (.A(_10224_),
    .B(_10217_),
    .Y(_10827_));
 sky130_fd_sc_hd__nor2_8 _33386_ (.A(_10223_),
    .B(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__a21o_2 _33387_ (.A1(_10821_),
    .A2(_10826_),
    .B1(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__nand3_4 _33388_ (.A(_10821_),
    .B(_10826_),
    .C(_10828_),
    .Y(_10830_));
 sky130_fd_sc_hd__nand2_1 _33389_ (.A(_10365_),
    .B(_10363_),
    .Y(_10831_));
 sky130_fd_sc_hd__nand2_4 _33390_ (.A(_10831_),
    .B(_10362_),
    .Y(_10832_));
 sky130_fd_sc_hd__a21oi_4 _33391_ (.A1(_10829_),
    .A2(_10830_),
    .B1(_10832_),
    .Y(_10833_));
 sky130_vsdinv _33392_ (.A(_10826_),
    .Y(_10834_));
 sky130_fd_sc_hd__nand2_2 _33393_ (.A(_10821_),
    .B(_10828_),
    .Y(_10835_));
 sky130_fd_sc_hd__o211a_2 _33394_ (.A1(_10834_),
    .A2(_10835_),
    .B1(_10832_),
    .C1(_10829_),
    .X(_10836_));
 sky130_fd_sc_hd__and2_4 _33395_ (.A(_10241_),
    .B(_10230_),
    .X(_10837_));
 sky130_fd_sc_hd__o21ai_4 _33396_ (.A1(_10833_),
    .A2(_10836_),
    .B1(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__nand2_1 _33397_ (.A(_10829_),
    .B(_10830_),
    .Y(_10839_));
 sky130_fd_sc_hd__and2_1 _33398_ (.A(_10831_),
    .B(_10362_),
    .X(_10840_));
 sky130_fd_sc_hd__nand2_1 _33399_ (.A(_10839_),
    .B(_10840_),
    .Y(_10841_));
 sky130_fd_sc_hd__nand3_4 _33400_ (.A(_10829_),
    .B(_10832_),
    .C(_10830_),
    .Y(_10842_));
 sky130_fd_sc_hd__nand3b_4 _33401_ (.A_N(_10837_),
    .B(_10841_),
    .C(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__o21ai_2 _33402_ (.A1(_10245_),
    .A2(_10239_),
    .B1(_10249_),
    .Y(_10844_));
 sky130_fd_sc_hd__a21oi_2 _33403_ (.A1(_10838_),
    .A2(_10843_),
    .B1(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__a21oi_1 _33404_ (.A1(_10246_),
    .A2(_10247_),
    .B1(_10245_),
    .Y(_10846_));
 sky130_fd_sc_hd__o211a_1 _33405_ (.A1(_10242_),
    .A2(_10846_),
    .B1(_10843_),
    .C1(_10838_),
    .X(_10847_));
 sky130_fd_sc_hd__o22ai_4 _33406_ (.A1(_10807_),
    .A2(_10808_),
    .B1(_10845_),
    .B2(_10847_),
    .Y(_10848_));
 sky130_fd_sc_hd__a21o_1 _33407_ (.A1(_10838_),
    .A2(_10843_),
    .B1(_10844_),
    .X(_10849_));
 sky130_fd_sc_hd__nor2_4 _33408_ (.A(_10807_),
    .B(_10808_),
    .Y(_10850_));
 sky130_fd_sc_hd__nand3_2 _33409_ (.A(_10838_),
    .B(_10844_),
    .C(_10843_),
    .Y(_10851_));
 sky130_fd_sc_hd__nand3_4 _33410_ (.A(_10849_),
    .B(_10850_),
    .C(_10851_),
    .Y(_10852_));
 sky130_fd_sc_hd__o21ai_4 _33411_ (.A1(_10378_),
    .A2(_10375_),
    .B1(_10376_),
    .Y(_10853_));
 sky130_fd_sc_hd__a21o_2 _33412_ (.A1(_10848_),
    .A2(_10852_),
    .B1(_10853_),
    .X(_10854_));
 sky130_fd_sc_hd__nand3_4 _33413_ (.A(_10848_),
    .B(_10853_),
    .C(_10852_),
    .Y(_10855_));
 sky130_fd_sc_hd__nand2_1 _33414_ (.A(_10298_),
    .B(_10292_),
    .Y(_10856_));
 sky130_fd_sc_hd__nand2_2 _33415_ (.A(_10856_),
    .B(_10297_),
    .Y(_10857_));
 sky130_fd_sc_hd__a21oi_1 _33416_ (.A1(_10854_),
    .A2(_10855_),
    .B1(_10857_),
    .Y(_10858_));
 sky130_fd_sc_hd__nand3_4 _33417_ (.A(_10854_),
    .B(_10855_),
    .C(_10857_),
    .Y(_10859_));
 sky130_vsdinv _33418_ (.A(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__o2bb2ai_2 _33419_ (.A1_N(_10751_),
    .A2_N(_10758_),
    .B1(_10858_),
    .B2(_10860_),
    .Y(_10861_));
 sky130_fd_sc_hd__nand2_1 _33420_ (.A(_10368_),
    .B(_10373_),
    .Y(_10862_));
 sky130_fd_sc_hd__a21oi_1 _33421_ (.A1(_10862_),
    .A2(_10488_),
    .B1(_10378_),
    .Y(_10863_));
 sky130_fd_sc_hd__o211a_2 _33422_ (.A1(_10491_),
    .A2(_10863_),
    .B1(_10852_),
    .C1(_10848_),
    .X(_10864_));
 sky130_fd_sc_hd__nand2_1 _33423_ (.A(_10854_),
    .B(_10857_),
    .Y(_10865_));
 sky130_fd_sc_hd__nor2_2 _33424_ (.A(_10254_),
    .B(_10292_),
    .Y(_10866_));
 sky130_fd_sc_hd__a21oi_4 _33425_ (.A1(_10848_),
    .A2(_10852_),
    .B1(_10853_),
    .Y(_10867_));
 sky130_fd_sc_hd__o22ai_4 _33426_ (.A1(_10251_),
    .A2(_10866_),
    .B1(_10867_),
    .B2(_10864_),
    .Y(_10868_));
 sky130_fd_sc_hd__o2111ai_4 _33427_ (.A1(_10864_),
    .A2(_10865_),
    .B1(_10868_),
    .C1(_10751_),
    .D1(_10758_),
    .Y(_10869_));
 sky130_fd_sc_hd__nand3_1 _33428_ (.A(_10306_),
    .B(_10500_),
    .C(_10308_),
    .Y(_10870_));
 sky130_fd_sc_hd__nand2_1 _33429_ (.A(_10870_),
    .B(_10511_),
    .Y(_10871_));
 sky130_fd_sc_hd__nand3_4 _33430_ (.A(_10861_),
    .B(_10869_),
    .C(_10871_),
    .Y(_10872_));
 sky130_fd_sc_hd__and2_1 _33431_ (.A(_10856_),
    .B(_10297_),
    .X(_10873_));
 sky130_fd_sc_hd__a21oi_2 _33432_ (.A1(_10854_),
    .A2(_10855_),
    .B1(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__nand2_2 _33433_ (.A(_10873_),
    .B(_10855_),
    .Y(_10875_));
 sky130_fd_sc_hd__nor2_2 _33434_ (.A(_10867_),
    .B(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__a21oi_4 _33435_ (.A1(_10745_),
    .A2(_10750_),
    .B1(_10747_),
    .Y(_10877_));
 sky130_fd_sc_hd__o211a_2 _33436_ (.A1(_10753_),
    .A2(_10754_),
    .B1(_10747_),
    .C1(_10745_),
    .X(_10878_));
 sky130_fd_sc_hd__o22ai_4 _33437_ (.A1(_10874_),
    .A2(_10876_),
    .B1(_10877_),
    .B2(_10878_),
    .Y(_10879_));
 sky130_fd_sc_hd__and3_1 _33438_ (.A(_10502_),
    .B(_10506_),
    .C(_10510_),
    .X(_10880_));
 sky130_fd_sc_hd__a31oi_4 _33439_ (.A1(_10308_),
    .A2(_10306_),
    .A3(_10500_),
    .B1(_10880_),
    .Y(_10881_));
 sky130_fd_sc_hd__nand2_2 _33440_ (.A(_10868_),
    .B(_10859_),
    .Y(_10882_));
 sky130_fd_sc_hd__nand3_2 _33441_ (.A(_10882_),
    .B(_10758_),
    .C(_10751_),
    .Y(_10883_));
 sky130_fd_sc_hd__nand3_4 _33442_ (.A(_10879_),
    .B(_10881_),
    .C(_10883_),
    .Y(_10884_));
 sky130_vsdinv _33443_ (.A(_10285_),
    .Y(_10885_));
 sky130_fd_sc_hd__nor2_8 _33444_ (.A(_10289_),
    .B(_10885_),
    .Y(_10886_));
 sky130_vsdinv _33445_ (.A(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__and2_2 _33446_ (.A(_10514_),
    .B(_10307_),
    .X(_10888_));
 sky130_fd_sc_hd__nor2_1 _33447_ (.A(_10887_),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__nand2_2 _33448_ (.A(_10514_),
    .B(_10307_),
    .Y(_10890_));
 sky130_fd_sc_hd__nor2_1 _33449_ (.A(_10886_),
    .B(_10890_),
    .Y(_10891_));
 sky130_fd_sc_hd__o2bb2ai_2 _33450_ (.A1_N(_10872_),
    .A2_N(_10884_),
    .B1(_10889_),
    .B2(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__a21boi_2 _33451_ (.A1(_10525_),
    .A2(_10209_),
    .B1_N(_10517_),
    .Y(_10893_));
 sky130_fd_sc_hd__nor2_4 _33452_ (.A(_10887_),
    .B(_10890_),
    .Y(_10894_));
 sky130_fd_sc_hd__nor2_8 _33453_ (.A(_10886_),
    .B(_10888_),
    .Y(_10895_));
 sky130_fd_sc_hd__nor2_4 _33454_ (.A(_10894_),
    .B(_10895_),
    .Y(_10896_));
 sky130_fd_sc_hd__nand3b_4 _33455_ (.A_N(_10896_),
    .B(_10884_),
    .C(_10872_),
    .Y(_10897_));
 sky130_fd_sc_hd__nand3_4 _33456_ (.A(_10892_),
    .B(_10893_),
    .C(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__o2bb2ai_2 _33457_ (.A1_N(_10872_),
    .A2_N(_10884_),
    .B1(_10895_),
    .B2(_10894_),
    .Y(_10899_));
 sky130_vsdinv _33458_ (.A(_10513_),
    .Y(_10900_));
 sky130_fd_sc_hd__nand2_1 _33459_ (.A(_10211_),
    .B(_10516_),
    .Y(_10901_));
 sky130_fd_sc_hd__o2bb2ai_2 _33460_ (.A1_N(_10525_),
    .A2_N(_10209_),
    .B1(_10900_),
    .B2(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__nand3_2 _33461_ (.A(_10884_),
    .B(_10872_),
    .C(_10896_),
    .Y(_10903_));
 sky130_fd_sc_hd__nand3_4 _33462_ (.A(_10899_),
    .B(_10902_),
    .C(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__nand3_2 _33463_ (.A(_10898_),
    .B(_10904_),
    .C(_10534_),
    .Y(_10905_));
 sky130_vsdinv _33464_ (.A(_10905_),
    .Y(_10906_));
 sky130_fd_sc_hd__o2bb2ai_2 _33465_ (.A1_N(_10904_),
    .A2_N(_10898_),
    .B1(_10529_),
    .B2(_10527_),
    .Y(_10907_));
 sky130_vsdinv _33466_ (.A(_10533_),
    .Y(_10908_));
 sky130_fd_sc_hd__o21ai_1 _33467_ (.A1(_10205_),
    .A2(_10175_),
    .B1(_10536_),
    .Y(_10909_));
 sky130_fd_sc_hd__o2bb2ai_2 _33468_ (.A1_N(_10538_),
    .A2_N(_10532_),
    .B1(_10908_),
    .B2(_10909_),
    .Y(_10910_));
 sky130_fd_sc_hd__nand2_4 _33469_ (.A(_10907_),
    .B(_10910_),
    .Y(_10911_));
 sky130_fd_sc_hd__a21o_2 _33470_ (.A1(_10907_),
    .A2(_10905_),
    .B1(_10910_),
    .X(_10912_));
 sky130_fd_sc_hd__o21ai_1 _33471_ (.A1(_10906_),
    .A2(_10911_),
    .B1(_10912_),
    .Y(_10913_));
 sky130_fd_sc_hd__and2b_1 _33472_ (.A_N(_10550_),
    .B(_10548_),
    .X(_10914_));
 sky130_fd_sc_hd__xor2_1 _33473_ (.A(_10913_),
    .B(_10914_),
    .X(_02650_));
 sky130_fd_sc_hd__o21a_4 _33474_ (.A1(_10753_),
    .A2(_10744_),
    .B1(_10666_),
    .X(_10915_));
 sky130_fd_sc_hd__buf_4 _33475_ (.A(_19857_),
    .X(_10916_));
 sky130_fd_sc_hd__buf_4 _33476_ (.A(_10916_),
    .X(_10917_));
 sky130_fd_sc_hd__buf_8 _33477_ (.A(_08775_),
    .X(_10918_));
 sky130_fd_sc_hd__clkbuf_4 _33478_ (.A(_06841_),
    .X(_10919_));
 sky130_fd_sc_hd__a22oi_4 _33479_ (.A1(_10917_),
    .A2(net454),
    .B1(_10918_),
    .B2(_10919_),
    .Y(_10920_));
 sky130_fd_sc_hd__nor2_4 _33480_ (.A(_06288_),
    .B(_10613_),
    .Y(_10921_));
 sky130_fd_sc_hd__nand2_4 _33481_ (.A(_07967_),
    .B(_06154_),
    .Y(_10922_));
 sky130_vsdinv _33482_ (.A(_10922_),
    .Y(_10923_));
 sky130_fd_sc_hd__o21ai_2 _33483_ (.A1(_10920_),
    .A2(_10921_),
    .B1(_10923_),
    .Y(_10924_));
 sky130_fd_sc_hd__a21oi_2 _33484_ (.A1(_10621_),
    .A2(_10616_),
    .B1(_10614_),
    .Y(_10925_));
 sky130_fd_sc_hd__buf_6 _33485_ (.A(_08775_),
    .X(_10926_));
 sky130_fd_sc_hd__a22o_2 _33486_ (.A1(_10917_),
    .A2(_06148_),
    .B1(_10926_),
    .B2(_10919_),
    .X(_10927_));
 sky130_fd_sc_hd__o211ai_2 _33487_ (.A1(_06298_),
    .A2(_10619_),
    .B1(_10922_),
    .C1(_10927_),
    .Y(_10928_));
 sky130_fd_sc_hd__nand3_4 _33488_ (.A(_10924_),
    .B(_10925_),
    .C(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__o21ai_2 _33489_ (.A1(_10920_),
    .A2(_10921_),
    .B1(_10922_),
    .Y(_10930_));
 sky130_fd_sc_hd__o211ai_2 _33490_ (.A1(_06298_),
    .A2(_10619_),
    .B1(_10923_),
    .C1(_10927_),
    .Y(_10931_));
 sky130_fd_sc_hd__o22ai_4 _33491_ (.A1(_10446_),
    .A2(_10619_),
    .B1(_10615_),
    .B2(_10612_),
    .Y(_10932_));
 sky130_fd_sc_hd__nand3_4 _33492_ (.A(_10930_),
    .B(_10931_),
    .C(_10932_),
    .Y(_10933_));
 sky130_fd_sc_hd__buf_4 _33493_ (.A(_19869_),
    .X(_10934_));
 sky130_fd_sc_hd__buf_6 _33494_ (.A(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__buf_4 _33495_ (.A(_08248_),
    .X(_10936_));
 sky130_fd_sc_hd__a22oi_4 _33496_ (.A1(_10935_),
    .A2(_20139_),
    .B1(_10936_),
    .B2(_20136_),
    .Y(_10937_));
 sky130_fd_sc_hd__nand2_2 _33497_ (.A(_10934_),
    .B(_07185_),
    .Y(_10938_));
 sky130_fd_sc_hd__nand2_2 _33498_ (.A(_19874_),
    .B(_06312_),
    .Y(_10939_));
 sky130_fd_sc_hd__nor2_2 _33499_ (.A(_10938_),
    .B(_10939_),
    .Y(_10940_));
 sky130_fd_sc_hd__buf_6 _33500_ (.A(_06715_),
    .X(_10941_));
 sky130_fd_sc_hd__nand2_2 _33501_ (.A(_07479_),
    .B(_10941_),
    .Y(_10942_));
 sky130_fd_sc_hd__o21bai_4 _33502_ (.A1(_10937_),
    .A2(_10940_),
    .B1_N(_10942_),
    .Y(_10943_));
 sky130_fd_sc_hd__buf_6 _33503_ (.A(_19872_),
    .X(_10944_));
 sky130_fd_sc_hd__buf_6 _33504_ (.A(_10944_),
    .X(_10945_));
 sky130_fd_sc_hd__nand3b_4 _33505_ (.A_N(_10938_),
    .B(_10945_),
    .C(_20136_),
    .Y(_10946_));
 sky130_fd_sc_hd__nand2_2 _33506_ (.A(_10938_),
    .B(_10939_),
    .Y(_10947_));
 sky130_fd_sc_hd__nand3_4 _33507_ (.A(_10946_),
    .B(_10942_),
    .C(_10947_),
    .Y(_10948_));
 sky130_fd_sc_hd__nand2_2 _33508_ (.A(_10943_),
    .B(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__a21o_2 _33509_ (.A1(_10929_),
    .A2(_10933_),
    .B1(_10949_),
    .X(_10950_));
 sky130_fd_sc_hd__nand3_4 _33510_ (.A(_10929_),
    .B(_10933_),
    .C(_10949_),
    .Y(_10951_));
 sky130_fd_sc_hd__nand2_4 _33511_ (.A(_10572_),
    .B(_10599_),
    .Y(_10952_));
 sky130_fd_sc_hd__a21o_2 _33512_ (.A1(_10950_),
    .A2(_10951_),
    .B1(_10952_),
    .X(_10953_));
 sky130_fd_sc_hd__nand3_4 _33513_ (.A(_10950_),
    .B(_10952_),
    .C(_10951_),
    .Y(_10954_));
 sky130_fd_sc_hd__a21boi_4 _33514_ (.A1(_10638_),
    .A2(_10623_),
    .B1_N(_10627_),
    .Y(_10955_));
 sky130_vsdinv _33515_ (.A(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__a21oi_2 _33516_ (.A1(_10953_),
    .A2(_10954_),
    .B1(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__and3_2 _33517_ (.A(_10950_),
    .B(_10952_),
    .C(_10951_),
    .X(_10958_));
 sky130_fd_sc_hd__nand2_2 _33518_ (.A(_10953_),
    .B(_10956_),
    .Y(_10959_));
 sky130_fd_sc_hd__nor2_2 _33519_ (.A(_10958_),
    .B(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__buf_4 _33520_ (.A(\pcpi_mul.rs2[32] ),
    .X(_10961_));
 sky130_fd_sc_hd__buf_4 _33521_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10962_));
 sky130_fd_sc_hd__nand3_4 _33522_ (.A(_10961_),
    .B(_10962_),
    .C(_05131_),
    .Y(_10963_));
 sky130_fd_sc_hd__nor2_2 _33523_ (.A(_05230_),
    .B(_10963_),
    .Y(_10964_));
 sky130_fd_sc_hd__nand2_4 _33524_ (.A(_10577_),
    .B(_05313_),
    .Y(_10965_));
 sky130_vsdinv _33525_ (.A(_10965_),
    .Y(_10966_));
 sky130_fd_sc_hd__clkinv_4 _33526_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_10967_));
 sky130_fd_sc_hd__buf_6 _33527_ (.A(_10967_),
    .X(_10968_));
 sky130_fd_sc_hd__o2bb2ai_4 _33528_ (.A1_N(_19829_),
    .A2_N(_20174_),
    .B1(_20177_),
    .B2(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__nand3b_1 _33529_ (.A_N(_10964_),
    .B(_10966_),
    .C(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__nand2_2 _33530_ (.A(_10970_),
    .B(_10579_),
    .Y(_10971_));
 sky130_fd_sc_hd__buf_6 _33531_ (.A(_10962_),
    .X(_10972_));
 sky130_fd_sc_hd__clkbuf_8 _33532_ (.A(_10961_),
    .X(_10973_));
 sky130_fd_sc_hd__a22oi_4 _33533_ (.A1(_10972_),
    .A2(_07901_),
    .B1(_04839_),
    .B2(_10973_),
    .Y(_10974_));
 sky130_fd_sc_hd__o21ai_2 _33534_ (.A1(_10964_),
    .A2(_10974_),
    .B1(_10966_),
    .Y(_10975_));
 sky130_vsdinv _33535_ (.A(_10579_),
    .Y(_10976_));
 sky130_fd_sc_hd__o211ai_4 _33536_ (.A1(_20178_),
    .A2(_10963_),
    .B1(_10965_),
    .C1(_10969_),
    .Y(_10977_));
 sky130_fd_sc_hd__nand3_4 _33537_ (.A(_10975_),
    .B(_10976_),
    .C(_10977_),
    .Y(_10978_));
 sky130_fd_sc_hd__nand2_4 _33538_ (.A(_09696_),
    .B(_05392_),
    .Y(_10979_));
 sky130_vsdinv _33539_ (.A(_10979_),
    .Y(_10980_));
 sky130_fd_sc_hd__a22oi_4 _33540_ (.A1(_09996_),
    .A2(_05451_),
    .B1(_10000_),
    .B2(_05283_),
    .Y(_10981_));
 sky130_fd_sc_hd__nand2_1 _33541_ (.A(\pcpi_mul.rs2[29] ),
    .B(\pcpi_mul.rs2[28] ),
    .Y(_10982_));
 sky130_fd_sc_hd__buf_6 _33542_ (.A(_10982_),
    .X(_10983_));
 sky130_fd_sc_hd__nor2_2 _33543_ (.A(_05862_),
    .B(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__nor2_1 _33544_ (.A(_10981_),
    .B(_10984_),
    .Y(_10985_));
 sky130_fd_sc_hd__nor2_1 _33545_ (.A(_10980_),
    .B(_10985_),
    .Y(_10986_));
 sky130_fd_sc_hd__buf_4 _33546_ (.A(_10982_),
    .X(_10987_));
 sky130_fd_sc_hd__buf_6 _33547_ (.A(_10987_),
    .X(_10988_));
 sky130_fd_sc_hd__buf_6 _33548_ (.A(_19839_),
    .X(_10989_));
 sky130_fd_sc_hd__a22o_2 _33549_ (.A1(_19835_),
    .A2(_05451_),
    .B1(_10989_),
    .B2(_05244_),
    .X(_10990_));
 sky130_fd_sc_hd__o211a_1 _33550_ (.A1(_05863_),
    .A2(_10988_),
    .B1(_10980_),
    .C1(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__o2bb2ai_2 _33551_ (.A1_N(_10971_),
    .A2_N(_10978_),
    .B1(_10986_),
    .B2(_10991_),
    .Y(_10992_));
 sky130_vsdinv _33552_ (.A(_10595_),
    .Y(_10993_));
 sky130_fd_sc_hd__o21ai_2 _33553_ (.A1(_10981_),
    .A2(_10984_),
    .B1(_10980_),
    .Y(_10994_));
 sky130_fd_sc_hd__o211ai_4 _33554_ (.A1(_05863_),
    .A2(_10987_),
    .B1(_10979_),
    .C1(_10990_),
    .Y(_10995_));
 sky130_fd_sc_hd__nand2_4 _33555_ (.A(_10994_),
    .B(_10995_),
    .Y(_10996_));
 sky130_fd_sc_hd__nand3_4 _33556_ (.A(_10978_),
    .B(_10971_),
    .C(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__nand3_4 _33557_ (.A(_10992_),
    .B(_10993_),
    .C(_10997_),
    .Y(_10998_));
 sky130_vsdinv _33558_ (.A(_10994_),
    .Y(_10999_));
 sky130_vsdinv _33559_ (.A(_10995_),
    .Y(_11000_));
 sky130_fd_sc_hd__o2bb2ai_1 _33560_ (.A1_N(_10971_),
    .A2_N(_10978_),
    .B1(_10999_),
    .B2(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__nand3b_1 _33561_ (.A_N(_10996_),
    .B(_10978_),
    .C(_10971_),
    .Y(_11002_));
 sky130_fd_sc_hd__nand3_2 _33562_ (.A(_11001_),
    .B(_10595_),
    .C(_11002_),
    .Y(_11003_));
 sky130_fd_sc_hd__buf_4 _33563_ (.A(_11003_),
    .X(_11004_));
 sky130_fd_sc_hd__or2_1 _33564_ (.A(_10561_),
    .B(_10556_),
    .X(_11005_));
 sky130_fd_sc_hd__nand2_1 _33565_ (.A(_08800_),
    .B(_05799_),
    .Y(_11006_));
 sky130_fd_sc_hd__nand3_2 _33566_ (.A(_11006_),
    .B(_10552_),
    .C(_05675_),
    .Y(_11007_));
 sky130_fd_sc_hd__buf_6 _33567_ (.A(_19846_),
    .X(_11008_));
 sky130_fd_sc_hd__nand2_1 _33568_ (.A(_11008_),
    .B(_06249_),
    .Y(_11009_));
 sky130_fd_sc_hd__buf_6 _33569_ (.A(_19850_),
    .X(_11010_));
 sky130_fd_sc_hd__nand3_2 _33570_ (.A(_11009_),
    .B(_11010_),
    .C(_05697_),
    .Y(_11011_));
 sky130_fd_sc_hd__o211ai_4 _33571_ (.A1(_08614_),
    .A2(_08243_),
    .B1(_11007_),
    .C1(_11011_),
    .Y(_11012_));
 sky130_fd_sc_hd__nand3_2 _33572_ (.A(_10552_),
    .B(_10384_),
    .C(_05577_),
    .Y(_11013_));
 sky130_fd_sc_hd__and2_1 _33573_ (.A(_19853_),
    .B(_05698_),
    .X(_11014_));
 sky130_fd_sc_hd__nand2_1 _33574_ (.A(_11009_),
    .B(_11006_),
    .Y(_11015_));
 sky130_fd_sc_hd__o211ai_4 _33575_ (.A1(_06256_),
    .A2(_11013_),
    .B1(_11014_),
    .C1(_11015_),
    .Y(_11016_));
 sky130_fd_sc_hd__nand2_1 _33576_ (.A(_11012_),
    .B(_11016_),
    .Y(_11017_));
 sky130_fd_sc_hd__o21ai_2 _33577_ (.A1(_10580_),
    .A2(_10582_),
    .B1(_10584_),
    .Y(_11018_));
 sky130_fd_sc_hd__nand2_1 _33578_ (.A(_11018_),
    .B(_10583_),
    .Y(_11019_));
 sky130_fd_sc_hd__nand2_1 _33579_ (.A(_11017_),
    .B(_11019_),
    .Y(_11020_));
 sky130_fd_sc_hd__o211ai_4 _33580_ (.A1(_10587_),
    .A2(_10592_),
    .B1(_11016_),
    .C1(_11012_),
    .Y(_11021_));
 sky130_fd_sc_hd__a22oi_4 _33581_ (.A1(_11005_),
    .A2(_10562_),
    .B1(_11020_),
    .B2(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__a21oi_4 _33582_ (.A1(_10562_),
    .A2(_10561_),
    .B1(_10556_),
    .Y(_11023_));
 sky130_fd_sc_hd__a22oi_4 _33583_ (.A1(_10583_),
    .A2(_11018_),
    .B1(_11012_),
    .B2(_11016_),
    .Y(_11024_));
 sky130_fd_sc_hd__nor2_2 _33584_ (.A(_11023_),
    .B(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__and2_1 _33585_ (.A(_11025_),
    .B(_11021_),
    .X(_11026_));
 sky130_fd_sc_hd__o2bb2ai_4 _33586_ (.A1_N(_10998_),
    .A2_N(_11004_),
    .B1(_11022_),
    .B2(_11026_),
    .Y(_11027_));
 sky130_fd_sc_hd__a21oi_4 _33587_ (.A1(_11021_),
    .A2(_11025_),
    .B1(_11022_),
    .Y(_11028_));
 sky130_fd_sc_hd__nand3_4 _33588_ (.A(_11028_),
    .B(_10998_),
    .C(_11004_),
    .Y(_11029_));
 sky130_fd_sc_hd__o211ai_2 _33589_ (.A1(_10564_),
    .A2(_10572_),
    .B1(_10598_),
    .C1(_10600_),
    .Y(_11030_));
 sky130_fd_sc_hd__nand2_4 _33590_ (.A(_11030_),
    .B(_10596_),
    .Y(_11031_));
 sky130_fd_sc_hd__a21oi_4 _33591_ (.A1(_11027_),
    .A2(_11029_),
    .B1(_11031_),
    .Y(_11032_));
 sky130_vsdinv _33592_ (.A(_10997_),
    .Y(_11033_));
 sky130_fd_sc_hd__nand2_1 _33593_ (.A(_10975_),
    .B(_10977_),
    .Y(_11034_));
 sky130_vsdinv _33594_ (.A(_10574_),
    .Y(_11035_));
 sky130_fd_sc_hd__nand2_2 _33595_ (.A(_10589_),
    .B(_10585_),
    .Y(_11036_));
 sky130_fd_sc_hd__o2111ai_4 _33596_ (.A1(_10996_),
    .A2(_11034_),
    .B1(_11035_),
    .C1(_10976_),
    .D1(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__nor2_1 _33597_ (.A(_11033_),
    .B(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand2_1 _33598_ (.A(_11028_),
    .B(_11004_),
    .Y(_11039_));
 sky130_fd_sc_hd__o211a_2 _33599_ (.A1(_11038_),
    .A2(_11039_),
    .B1(_11031_),
    .C1(_11027_),
    .X(_11040_));
 sky130_fd_sc_hd__o22ai_4 _33600_ (.A1(_10957_),
    .A2(_10960_),
    .B1(_11032_),
    .B2(_11040_),
    .Y(_11041_));
 sky130_fd_sc_hd__a21oi_2 _33601_ (.A1(_10998_),
    .A2(_11004_),
    .B1(_11028_),
    .Y(_11042_));
 sky130_fd_sc_hd__o211a_1 _33602_ (.A1(_11033_),
    .A2(_11037_),
    .B1(_11028_),
    .C1(_11003_),
    .X(_11043_));
 sky130_fd_sc_hd__o21bai_4 _33603_ (.A1(_11042_),
    .A2(_11043_),
    .B1_N(_11031_),
    .Y(_11044_));
 sky130_fd_sc_hd__a21oi_4 _33604_ (.A1(_10950_),
    .A2(_10951_),
    .B1(_10952_),
    .Y(_11045_));
 sky130_fd_sc_hd__o21ai_2 _33605_ (.A1(_11045_),
    .A2(_10958_),
    .B1(_10956_),
    .Y(_11046_));
 sky130_fd_sc_hd__nand3_2 _33606_ (.A(_10953_),
    .B(_10954_),
    .C(_10955_),
    .Y(_11047_));
 sky130_fd_sc_hd__nand2_4 _33607_ (.A(_11046_),
    .B(_11047_),
    .Y(_11048_));
 sky130_fd_sc_hd__nand3_4 _33608_ (.A(_11027_),
    .B(_11029_),
    .C(_11031_),
    .Y(_11049_));
 sky130_fd_sc_hd__nand3_4 _33609_ (.A(_11044_),
    .B(_11048_),
    .C(_11049_),
    .Y(_11050_));
 sky130_fd_sc_hd__nand2_4 _33610_ (.A(_10660_),
    .B(_10606_),
    .Y(_11051_));
 sky130_fd_sc_hd__a21oi_4 _33611_ (.A1(_11041_),
    .A2(_11050_),
    .B1(_11051_),
    .Y(_11052_));
 sky130_fd_sc_hd__nand2_1 _33612_ (.A(_11044_),
    .B(_11048_),
    .Y(_11053_));
 sky130_fd_sc_hd__o211a_1 _33613_ (.A1(_11040_),
    .A2(_11053_),
    .B1(_11051_),
    .C1(_11041_),
    .X(_11054_));
 sky130_fd_sc_hd__nor2_1 _33614_ (.A(_10725_),
    .B(_10687_),
    .Y(_11055_));
 sky130_fd_sc_hd__a21oi_2 _33615_ (.A1(_10652_),
    .A2(_10655_),
    .B1(_10645_),
    .Y(_11056_));
 sky130_fd_sc_hd__buf_6 _33616_ (.A(_09602_),
    .X(_11057_));
 sky130_fd_sc_hd__clkbuf_4 _33617_ (.A(_06543_),
    .X(_11058_));
 sky130_fd_sc_hd__nand3_4 _33618_ (.A(_11058_),
    .B(_07422_),
    .C(_07250_),
    .Y(_11059_));
 sky130_fd_sc_hd__nor2_8 _33619_ (.A(_11057_),
    .B(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__clkbuf_4 _33620_ (.A(_07254_),
    .X(_11061_));
 sky130_fd_sc_hd__clkbuf_4 _33621_ (.A(_20114_),
    .X(_11062_));
 sky130_fd_sc_hd__a22o_2 _33622_ (.A1(_06358_),
    .A2(_11061_),
    .B1(_10693_),
    .B2(_11062_),
    .X(_11063_));
 sky130_fd_sc_hd__nand2_2 _33623_ (.A(_10700_),
    .B(_08056_),
    .Y(_11064_));
 sky130_vsdinv _33624_ (.A(_11064_),
    .Y(_11065_));
 sky130_fd_sc_hd__nand2_1 _33625_ (.A(_11063_),
    .B(_11065_),
    .Y(_11066_));
 sky130_fd_sc_hd__a22oi_4 _33626_ (.A1(_06358_),
    .A2(_20119_),
    .B1(_10351_),
    .B2(_11062_),
    .Y(_11067_));
 sky130_fd_sc_hd__o21ai_2 _33627_ (.A1(_11067_),
    .A2(_11060_),
    .B1(_11064_),
    .Y(_11068_));
 sky130_fd_sc_hd__nor2_2 _33628_ (.A(_10696_),
    .B(_10697_),
    .Y(_11069_));
 sky130_fd_sc_hd__a21o_1 _33629_ (.A1(_10702_),
    .A2(_10698_),
    .B1(_11069_),
    .X(_11070_));
 sky130_fd_sc_hd__o211ai_4 _33630_ (.A1(_11060_),
    .A2(_11066_),
    .B1(_11068_),
    .C1(_11070_),
    .Y(_11071_));
 sky130_fd_sc_hd__o21ai_2 _33631_ (.A1(_11067_),
    .A2(_11060_),
    .B1(_11065_),
    .Y(_11072_));
 sky130_fd_sc_hd__a21oi_2 _33632_ (.A1(_10702_),
    .A2(_10698_),
    .B1(_11069_),
    .Y(_11073_));
 sky130_fd_sc_hd__buf_6 _33633_ (.A(_11057_),
    .X(_11074_));
 sky130_fd_sc_hd__o211ai_4 _33634_ (.A1(_11074_),
    .A2(_11059_),
    .B1(_11064_),
    .C1(_11063_),
    .Y(_11075_));
 sky130_fd_sc_hd__nand3_4 _33635_ (.A(_11072_),
    .B(_11073_),
    .C(_11075_),
    .Y(_11076_));
 sky130_fd_sc_hd__nand2_1 _33636_ (.A(_11071_),
    .B(_11076_),
    .Y(_11077_));
 sky130_fd_sc_hd__buf_6 _33637_ (.A(_08450_),
    .X(_11078_));
 sky130_fd_sc_hd__a22oi_4 _33638_ (.A1(_10337_),
    .A2(_20108_),
    .B1(_10338_),
    .B2(_11078_),
    .Y(_11079_));
 sky130_fd_sc_hd__nand2_2 _33639_ (.A(_06531_),
    .B(_08052_),
    .Y(_11080_));
 sky130_fd_sc_hd__nand2_1 _33640_ (.A(_19906_),
    .B(_10716_),
    .Y(_11081_));
 sky130_fd_sc_hd__nor2_1 _33641_ (.A(_11080_),
    .B(_11081_),
    .Y(_11082_));
 sky130_fd_sc_hd__nand2_2 _33642_ (.A(_05953_),
    .B(_10811_),
    .Y(_11083_));
 sky130_fd_sc_hd__o21bai_2 _33643_ (.A1(_11079_),
    .A2(_11082_),
    .B1_N(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__buf_4 _33644_ (.A(_09926_),
    .X(_11085_));
 sky130_fd_sc_hd__nand3b_4 _33645_ (.A_N(_11080_),
    .B(_19907_),
    .C(_11085_),
    .Y(_11086_));
 sky130_fd_sc_hd__nand2_1 _33646_ (.A(_11080_),
    .B(_11081_),
    .Y(_11087_));
 sky130_fd_sc_hd__nand3_2 _33647_ (.A(_11086_),
    .B(_11083_),
    .C(_11087_),
    .Y(_11088_));
 sky130_fd_sc_hd__nand2_4 _33648_ (.A(_11084_),
    .B(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__and2_1 _33649_ (.A(_11077_),
    .B(_11089_),
    .X(_11090_));
 sky130_fd_sc_hd__nor2_2 _33650_ (.A(_11089_),
    .B(_11077_),
    .Y(_11091_));
 sky130_fd_sc_hd__buf_6 _33651_ (.A(_07754_),
    .X(_11092_));
 sky130_fd_sc_hd__buf_4 _33652_ (.A(_06719_),
    .X(_11093_));
 sky130_fd_sc_hd__buf_6 _33653_ (.A(_06637_),
    .X(_11094_));
 sky130_fd_sc_hd__a22oi_4 _33654_ (.A1(_11092_),
    .A2(_11093_),
    .B1(_11094_),
    .B2(_07258_),
    .Y(_11095_));
 sky130_vsdinv _33655_ (.A(_08142_),
    .Y(_11096_));
 sky130_fd_sc_hd__nor2_4 _33656_ (.A(_11096_),
    .B(_10668_),
    .Y(_11097_));
 sky130_fd_sc_hd__nand2_2 _33657_ (.A(_19890_),
    .B(_07567_),
    .Y(_11098_));
 sky130_vsdinv _33658_ (.A(_11098_),
    .Y(_11099_));
 sky130_fd_sc_hd__o21ai_2 _33659_ (.A1(_11095_),
    .A2(_11097_),
    .B1(_11099_),
    .Y(_11100_));
 sky130_fd_sc_hd__nand2_1 _33660_ (.A(_10630_),
    .B(_10631_),
    .Y(_11101_));
 sky130_fd_sc_hd__a21oi_4 _33661_ (.A1(_10636_),
    .A2(_11101_),
    .B1(_10632_),
    .Y(_11102_));
 sky130_fd_sc_hd__buf_4 _33662_ (.A(_07754_),
    .X(_11103_));
 sky130_fd_sc_hd__a22o_2 _33663_ (.A1(_11103_),
    .A2(_11093_),
    .B1(_11094_),
    .B2(_07258_),
    .X(_11104_));
 sky130_fd_sc_hd__o211ai_4 _33664_ (.A1(_11096_),
    .A2(_10668_),
    .B1(_11098_),
    .C1(_11104_),
    .Y(_11105_));
 sky130_fd_sc_hd__nand3_4 _33665_ (.A(_11100_),
    .B(_11102_),
    .C(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__o21ai_2 _33666_ (.A1(_11095_),
    .A2(_11097_),
    .B1(_11098_),
    .Y(_11107_));
 sky130_fd_sc_hd__nand3b_1 _33667_ (.A_N(_10630_),
    .B(_10936_),
    .C(_20139_),
    .Y(_11108_));
 sky130_fd_sc_hd__o21ai_2 _33668_ (.A1(_10634_),
    .A2(_10629_),
    .B1(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__o211ai_4 _33669_ (.A1(_11096_),
    .A2(_10668_),
    .B1(_11099_),
    .C1(_11104_),
    .Y(_11110_));
 sky130_fd_sc_hd__nand3_4 _33670_ (.A(_11107_),
    .B(_11109_),
    .C(_11110_),
    .Y(_11111_));
 sky130_vsdinv _33671_ (.A(_10669_),
    .Y(_11112_));
 sky130_fd_sc_hd__nor2_4 _33672_ (.A(_10672_),
    .B(_10678_),
    .Y(_11113_));
 sky130_fd_sc_hd__o2bb2ai_4 _33673_ (.A1_N(_11106_),
    .A2_N(_11111_),
    .B1(_11112_),
    .B2(_11113_),
    .Y(_11114_));
 sky130_fd_sc_hd__nor2_2 _33674_ (.A(_11112_),
    .B(_11113_),
    .Y(_11115_));
 sky130_fd_sc_hd__nand3_4 _33675_ (.A(_11106_),
    .B(_11111_),
    .C(_11115_),
    .Y(_11116_));
 sky130_vsdinv _33676_ (.A(_10683_),
    .Y(_11117_));
 sky130_fd_sc_hd__nand2_1 _33677_ (.A(_10676_),
    .B(_11117_),
    .Y(_11118_));
 sky130_fd_sc_hd__nand2_4 _33678_ (.A(_11118_),
    .B(_10680_),
    .Y(_11119_));
 sky130_fd_sc_hd__a21oi_4 _33679_ (.A1(_11114_),
    .A2(_11116_),
    .B1(_11119_),
    .Y(_11120_));
 sky130_fd_sc_hd__a21oi_1 _33680_ (.A1(_10673_),
    .A2(_10675_),
    .B1(_10674_),
    .Y(_11121_));
 sky130_fd_sc_hd__o211a_1 _33681_ (.A1(_11121_),
    .A2(_10684_),
    .B1(_11116_),
    .C1(_11114_),
    .X(_11122_));
 sky130_fd_sc_hd__o22ai_4 _33682_ (.A1(_11090_),
    .A2(_11091_),
    .B1(_11120_),
    .B2(_11122_),
    .Y(_11123_));
 sky130_fd_sc_hd__a21o_1 _33683_ (.A1(_11114_),
    .A2(_11116_),
    .B1(_11119_),
    .X(_11124_));
 sky130_fd_sc_hd__nand3_4 _33684_ (.A(_11119_),
    .B(_11114_),
    .C(_11116_),
    .Y(_11125_));
 sky130_vsdinv _33685_ (.A(_11071_),
    .Y(_11126_));
 sky130_fd_sc_hd__nand2_2 _33686_ (.A(_11076_),
    .B(_11089_),
    .Y(_11127_));
 sky130_fd_sc_hd__a21o_1 _33687_ (.A1(_11071_),
    .A2(_11076_),
    .B1(_11089_),
    .X(_11128_));
 sky130_fd_sc_hd__o21ai_4 _33688_ (.A1(_11126_),
    .A2(_11127_),
    .B1(_11128_),
    .Y(_11129_));
 sky130_fd_sc_hd__nand3_4 _33689_ (.A(_11124_),
    .B(_11125_),
    .C(_11129_),
    .Y(_11130_));
 sky130_fd_sc_hd__nand3_4 _33690_ (.A(_11056_),
    .B(_11123_),
    .C(_11130_),
    .Y(_11131_));
 sky130_fd_sc_hd__o21a_2 _33691_ (.A1(_10690_),
    .A2(_11055_),
    .B1(_11131_),
    .X(_11132_));
 sky130_fd_sc_hd__o21ai_2 _33692_ (.A1(_11120_),
    .A2(_11122_),
    .B1(_11129_),
    .Y(_11133_));
 sky130_vsdinv _33693_ (.A(_10655_),
    .Y(_11134_));
 sky130_fd_sc_hd__o21ai_2 _33694_ (.A1(_11134_),
    .A2(_10643_),
    .B1(_10653_),
    .Y(_11135_));
 sky130_fd_sc_hd__nand3b_2 _33695_ (.A_N(_11129_),
    .B(_11124_),
    .C(_11125_),
    .Y(_11136_));
 sky130_fd_sc_hd__nand3_4 _33696_ (.A(_11133_),
    .B(_11135_),
    .C(_11136_),
    .Y(_11137_));
 sky130_fd_sc_hd__o21ai_4 _33697_ (.A1(_10725_),
    .A2(_10687_),
    .B1(_10731_),
    .Y(_11138_));
 sky130_fd_sc_hd__a21oi_4 _33698_ (.A1(_11137_),
    .A2(_11131_),
    .B1(_11138_),
    .Y(_11139_));
 sky130_fd_sc_hd__a21oi_4 _33699_ (.A1(_11132_),
    .A2(_11137_),
    .B1(_11139_),
    .Y(_11140_));
 sky130_fd_sc_hd__o21ai_2 _33700_ (.A1(_11052_),
    .A2(_11054_),
    .B1(_11140_),
    .Y(_11141_));
 sky130_fd_sc_hd__a21o_2 _33701_ (.A1(_11041_),
    .A2(_11050_),
    .B1(_11051_),
    .X(_11142_));
 sky130_fd_sc_hd__nand3_4 _33702_ (.A(_11041_),
    .B(_11051_),
    .C(_11050_),
    .Y(_11143_));
 sky130_fd_sc_hd__a22oi_4 _33703_ (.A1(_10656_),
    .A2(_10653_),
    .B1(_11123_),
    .B2(_11130_),
    .Y(_11144_));
 sky130_fd_sc_hd__nand2_2 _33704_ (.A(_11131_),
    .B(_11138_),
    .Y(_11145_));
 sky130_fd_sc_hd__a21o_1 _33705_ (.A1(_11137_),
    .A2(_11131_),
    .B1(_11138_),
    .X(_11146_));
 sky130_fd_sc_hd__o21ai_2 _33706_ (.A1(_11144_),
    .A2(_11145_),
    .B1(_11146_),
    .Y(_11147_));
 sky130_fd_sc_hd__nand3_2 _33707_ (.A(_11142_),
    .B(_11143_),
    .C(_11147_),
    .Y(_11148_));
 sky130_fd_sc_hd__nand3_4 _33708_ (.A(_10915_),
    .B(_11141_),
    .C(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__nor2_2 _33709_ (.A(_11144_),
    .B(_11145_),
    .Y(_11150_));
 sky130_fd_sc_hd__o22ai_4 _33710_ (.A1(_11150_),
    .A2(_11139_),
    .B1(_11052_),
    .B2(_11054_),
    .Y(_11151_));
 sky130_fd_sc_hd__o21ai_4 _33711_ (.A1(_10753_),
    .A2(_10744_),
    .B1(_10666_),
    .Y(_11152_));
 sky130_fd_sc_hd__nand3_4 _33712_ (.A(_11142_),
    .B(_11143_),
    .C(_11140_),
    .Y(_11153_));
 sky130_fd_sc_hd__nand3_2 _33713_ (.A(_11151_),
    .B(_11152_),
    .C(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__nand2_2 _33714_ (.A(_11149_),
    .B(_11154_),
    .Y(_11155_));
 sky130_fd_sc_hd__nand2_2 _33715_ (.A(_19921_),
    .B(_09787_),
    .Y(_11156_));
 sky130_fd_sc_hd__buf_6 _33716_ (.A(_20081_),
    .X(_11157_));
 sky130_fd_sc_hd__nand2_2 _33717_ (.A(_05805_),
    .B(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__nor2_2 _33718_ (.A(_11156_),
    .B(_11158_),
    .Y(_11159_));
 sky130_fd_sc_hd__nand2_4 _33719_ (.A(_18685_),
    .B(net469),
    .Y(_11160_));
 sky130_fd_sc_hd__inv_2 _33720_ (.A(_11160_),
    .Y(_11161_));
 sky130_fd_sc_hd__buf_2 _33721_ (.A(_11161_),
    .X(_11162_));
 sky130_fd_sc_hd__nand2_2 _33722_ (.A(_11156_),
    .B(_11158_),
    .Y(_11163_));
 sky130_fd_sc_hd__nand3b_4 _33723_ (.A_N(_11159_),
    .B(_11162_),
    .C(_11163_),
    .Y(_11164_));
 sky130_fd_sc_hd__buf_8 _33724_ (.A(_09896_),
    .X(_11165_));
 sky130_fd_sc_hd__a21o_1 _33725_ (.A1(_19926_),
    .A2(_11165_),
    .B1(_11156_),
    .X(_11166_));
 sky130_fd_sc_hd__a21o_1 _33726_ (.A1(_19921_),
    .A2(_20087_),
    .B1(_11158_),
    .X(_11167_));
 sky130_fd_sc_hd__clkbuf_4 _33727_ (.A(_11160_),
    .X(_11168_));
 sky130_fd_sc_hd__nand3_4 _33728_ (.A(_11166_),
    .B(_11167_),
    .C(_11168_),
    .Y(_11169_));
 sky130_fd_sc_hd__a21o_2 _33729_ (.A1(_10789_),
    .A2(_10785_),
    .B1(_10793_),
    .X(_11170_));
 sky130_fd_sc_hd__a21oi_4 _33730_ (.A1(_11164_),
    .A2(_11169_),
    .B1(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__and3_1 _33731_ (.A(_11164_),
    .B(_11170_),
    .C(_11169_),
    .X(_11172_));
 sky130_fd_sc_hd__buf_4 _33732_ (.A(\pcpi_mul.rs1[30] ),
    .X(_11173_));
 sky130_fd_sc_hd__buf_4 _33733_ (.A(_11173_),
    .X(_11174_));
 sky130_fd_sc_hd__and4_1 _33734_ (.A(_05140_),
    .B(_05142_),
    .C(_10778_),
    .D(_11174_),
    .X(_11175_));
 sky130_vsdinv _33735_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_11176_));
 sky130_fd_sc_hd__buf_6 _33736_ (.A(_11176_),
    .X(_11177_));
 sky130_fd_sc_hd__nand2_1 _33737_ (.A(_19932_),
    .B(_20074_),
    .Y(_11178_));
 sky130_fd_sc_hd__o21a_1 _33738_ (.A1(_05151_),
    .A2(_11177_),
    .B1(_11178_),
    .X(_11179_));
 sky130_vsdinv _33739_ (.A(\pcpi_mul.rs1[29] ),
    .Y(_11180_));
 sky130_fd_sc_hd__buf_8 _33740_ (.A(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__nor2_4 _33741_ (.A(_05154_),
    .B(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__o21bai_2 _33742_ (.A1(_11175_),
    .A2(_11179_),
    .B1_N(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__o21ai_2 _33743_ (.A1(_05151_),
    .A2(_11177_),
    .B1(_11178_),
    .Y(_11184_));
 sky130_fd_sc_hd__nand3b_4 _33744_ (.A_N(_11175_),
    .B(_11182_),
    .C(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__nand2_4 _33745_ (.A(_11183_),
    .B(_11185_),
    .Y(_11186_));
 sky130_fd_sc_hd__o21ai_4 _33746_ (.A1(_11171_),
    .A2(_11172_),
    .B1(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__nand2_1 _33747_ (.A(_10792_),
    .B(_10775_),
    .Y(_11188_));
 sky130_fd_sc_hd__nand2_2 _33748_ (.A(_11188_),
    .B(_10796_),
    .Y(_11189_));
 sky130_fd_sc_hd__and2_1 _33749_ (.A(_11183_),
    .B(_11185_),
    .X(_11190_));
 sky130_fd_sc_hd__a21o_1 _33750_ (.A1(_11164_),
    .A2(_11169_),
    .B1(_11170_),
    .X(_11191_));
 sky130_fd_sc_hd__nand3_4 _33751_ (.A(_11164_),
    .B(_11170_),
    .C(_11169_),
    .Y(_11192_));
 sky130_fd_sc_hd__nand3_4 _33752_ (.A(_11190_),
    .B(_11191_),
    .C(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__nand3_4 _33753_ (.A(_11187_),
    .B(_11189_),
    .C(_11193_),
    .Y(_11194_));
 sky130_fd_sc_hd__o21ai_2 _33754_ (.A1(_11171_),
    .A2(_11172_),
    .B1(_11190_),
    .Y(_11195_));
 sky130_fd_sc_hd__a21boi_4 _33755_ (.A1(_10792_),
    .A2(_10775_),
    .B1_N(_10796_),
    .Y(_11196_));
 sky130_fd_sc_hd__nand3_2 _33756_ (.A(_11191_),
    .B(_11192_),
    .C(_11186_),
    .Y(_11197_));
 sky130_fd_sc_hd__nand3_4 _33757_ (.A(_11195_),
    .B(_11196_),
    .C(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__a21oi_4 _33758_ (.A1(_10770_),
    .A2(_10764_),
    .B1(_10762_),
    .Y(_11199_));
 sky130_fd_sc_hd__a21boi_4 _33759_ (.A1(_11194_),
    .A2(_11198_),
    .B1_N(_11199_),
    .Y(_11200_));
 sky130_fd_sc_hd__a31oi_4 _33760_ (.A1(_11187_),
    .A2(_11189_),
    .A3(_11193_),
    .B1(_11199_),
    .Y(_11201_));
 sky130_fd_sc_hd__and2_2 _33761_ (.A(_11201_),
    .B(_11198_),
    .X(_11202_));
 sky130_vsdinv _33762_ (.A(_10821_),
    .Y(_11203_));
 sky130_fd_sc_hd__nor2_2 _33763_ (.A(_10828_),
    .B(_10834_),
    .Y(_11204_));
 sky130_fd_sc_hd__buf_4 _33764_ (.A(_20097_),
    .X(_11205_));
 sky130_fd_sc_hd__clkbuf_4 _33765_ (.A(_19915_),
    .X(_11206_));
 sky130_fd_sc_hd__a22oi_4 _33766_ (.A1(_10809_),
    .A2(_11205_),
    .B1(_11206_),
    .B2(_20094_),
    .Y(_11207_));
 sky130_fd_sc_hd__nand3_4 _33767_ (.A(_05858_),
    .B(_05608_),
    .C(_09490_),
    .Y(_11208_));
 sky130_fd_sc_hd__nor2_4 _33768_ (.A(_08888_),
    .B(_11208_),
    .Y(_11209_));
 sky130_fd_sc_hd__buf_6 _33769_ (.A(\pcpi_mul.rs1[26] ),
    .X(_11210_));
 sky130_fd_sc_hd__nand2_2 _33770_ (.A(_05866_),
    .B(_11210_),
    .Y(_11211_));
 sky130_fd_sc_hd__o21ai_2 _33771_ (.A1(_11207_),
    .A2(_11209_),
    .B1(_11211_),
    .Y(_11212_));
 sky130_vsdinv _33772_ (.A(_11211_),
    .Y(_11213_));
 sky130_fd_sc_hd__a22o_1 _33773_ (.A1(_19913_),
    .A2(_20098_),
    .B1(_11206_),
    .B2(_20094_),
    .X(_11214_));
 sky130_fd_sc_hd__o211ai_2 _33774_ (.A1(_08888_),
    .A2(_11208_),
    .B1(_11213_),
    .C1(_11214_),
    .Y(_11215_));
 sky130_fd_sc_hd__o21ai_2 _33775_ (.A1(_10717_),
    .A2(_10712_),
    .B1(_10719_),
    .Y(_11216_));
 sky130_fd_sc_hd__nand3_4 _33776_ (.A(_11212_),
    .B(_11215_),
    .C(_11216_),
    .Y(_11217_));
 sky130_fd_sc_hd__o21ai_2 _33777_ (.A1(_11207_),
    .A2(_11209_),
    .B1(_11213_),
    .Y(_11218_));
 sky130_fd_sc_hd__o21ai_1 _33778_ (.A1(_10713_),
    .A2(_10714_),
    .B1(_10717_),
    .Y(_11219_));
 sky130_fd_sc_hd__nand2_2 _33779_ (.A(_11219_),
    .B(_10720_),
    .Y(_11220_));
 sky130_fd_sc_hd__o211ai_2 _33780_ (.A1(_09880_),
    .A2(_11208_),
    .B1(_11211_),
    .C1(_11214_),
    .Y(_11221_));
 sky130_fd_sc_hd__nand3_4 _33781_ (.A(_11218_),
    .B(_11220_),
    .C(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__nor2_4 _33782_ (.A(_10816_),
    .B(_10813_),
    .Y(_11223_));
 sky130_fd_sc_hd__o2bb2ai_4 _33783_ (.A1_N(_11217_),
    .A2_N(_11222_),
    .B1(_10810_),
    .B2(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__nor2_2 _33784_ (.A(_10810_),
    .B(_11223_),
    .Y(_11225_));
 sky130_fd_sc_hd__nand3_4 _33785_ (.A(_11217_),
    .B(_11222_),
    .C(_11225_),
    .Y(_11226_));
 sky130_fd_sc_hd__nand2_4 _33786_ (.A(_10723_),
    .B(_10708_),
    .Y(_11227_));
 sky130_fd_sc_hd__a21oi_4 _33787_ (.A1(_11224_),
    .A2(_11226_),
    .B1(_11227_),
    .Y(_11228_));
 sky130_fd_sc_hd__nand2_1 _33788_ (.A(_11222_),
    .B(_11225_),
    .Y(_11229_));
 sky130_vsdinv _33789_ (.A(_11217_),
    .Y(_11230_));
 sky130_fd_sc_hd__o211a_2 _33790_ (.A1(_11229_),
    .A2(_11230_),
    .B1(_11224_),
    .C1(_11227_),
    .X(_11231_));
 sky130_fd_sc_hd__o22ai_4 _33791_ (.A1(_11203_),
    .A2(_11204_),
    .B1(_11228_),
    .B2(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__a21o_1 _33792_ (.A1(_11224_),
    .A2(_11226_),
    .B1(_11227_),
    .X(_11233_));
 sky130_fd_sc_hd__nand3_4 _33793_ (.A(_11227_),
    .B(_11224_),
    .C(_11226_),
    .Y(_11234_));
 sky130_fd_sc_hd__nand2_4 _33794_ (.A(_10835_),
    .B(_10826_),
    .Y(_11235_));
 sky130_fd_sc_hd__nand3_4 _33795_ (.A(_11233_),
    .B(_11234_),
    .C(_11235_),
    .Y(_11236_));
 sky130_fd_sc_hd__o21ai_4 _33796_ (.A1(_10837_),
    .A2(_10833_),
    .B1(_10842_),
    .Y(_11237_));
 sky130_fd_sc_hd__a21oi_4 _33797_ (.A1(_11232_),
    .A2(_11236_),
    .B1(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__a21oi_2 _33798_ (.A1(_10839_),
    .A2(_10840_),
    .B1(_10837_),
    .Y(_11239_));
 sky130_fd_sc_hd__o211a_4 _33799_ (.A1(_10836_),
    .A2(_11239_),
    .B1(_11236_),
    .C1(_11232_),
    .X(_11240_));
 sky130_fd_sc_hd__o22ai_4 _33800_ (.A1(_11200_),
    .A2(_11202_),
    .B1(_11238_),
    .B2(_11240_),
    .Y(_11241_));
 sky130_fd_sc_hd__a21o_1 _33801_ (.A1(_11232_),
    .A2(_11236_),
    .B1(_11237_),
    .X(_11242_));
 sky130_fd_sc_hd__a21oi_4 _33802_ (.A1(_11198_),
    .A2(_11201_),
    .B1(_11200_),
    .Y(_11243_));
 sky130_fd_sc_hd__nand3_4 _33803_ (.A(_11237_),
    .B(_11232_),
    .C(_11236_),
    .Y(_11244_));
 sky130_fd_sc_hd__nand3_4 _33804_ (.A(_11242_),
    .B(_11243_),
    .C(_11244_),
    .Y(_11245_));
 sky130_vsdinv _33805_ (.A(_10732_),
    .Y(_11246_));
 sky130_fd_sc_hd__nand2_1 _33806_ (.A(_10726_),
    .B(_10728_),
    .Y(_11247_));
 sky130_fd_sc_hd__o2bb2ai_4 _33807_ (.A1_N(_10740_),
    .A2_N(_10741_),
    .B1(_11246_),
    .B2(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__a21oi_4 _33808_ (.A1(_11241_),
    .A2(_11245_),
    .B1(_11248_),
    .Y(_11249_));
 sky130_fd_sc_hd__nand2_1 _33809_ (.A(_11243_),
    .B(_11244_),
    .Y(_11250_));
 sky130_fd_sc_hd__o211a_2 _33810_ (.A1(_11238_),
    .A2(_11250_),
    .B1(_11248_),
    .C1(_11241_),
    .X(_11251_));
 sky130_fd_sc_hd__a21o_4 _33811_ (.A1(_10849_),
    .A2(_10850_),
    .B1(_10847_),
    .X(_11252_));
 sky130_fd_sc_hd__o21bai_4 _33812_ (.A1(_11249_),
    .A2(_11251_),
    .B1_N(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__a21o_1 _33813_ (.A1(_11241_),
    .A2(_11245_),
    .B1(_11248_),
    .X(_11254_));
 sky130_fd_sc_hd__nand3_4 _33814_ (.A(_11241_),
    .B(_11248_),
    .C(_11245_),
    .Y(_11255_));
 sky130_fd_sc_hd__nand3_4 _33815_ (.A(_11254_),
    .B(_11255_),
    .C(_11252_),
    .Y(_11256_));
 sky130_fd_sc_hd__nand2_8 _33816_ (.A(_11253_),
    .B(_11256_),
    .Y(_11257_));
 sky130_fd_sc_hd__nand2_8 _33817_ (.A(_11155_),
    .B(_11257_),
    .Y(_11258_));
 sky130_fd_sc_hd__nand2_1 _33818_ (.A(_10747_),
    .B(_10750_),
    .Y(_11259_));
 sky130_fd_sc_hd__o22ai_4 _33819_ (.A1(_10752_),
    .A2(_11259_),
    .B1(_10877_),
    .B2(_10882_),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_2 _33820_ (.A(_11254_),
    .B(_11252_),
    .Y(_11261_));
 sky130_fd_sc_hd__buf_4 _33821_ (.A(_11154_),
    .X(_11262_));
 sky130_fd_sc_hd__o2111ai_4 _33822_ (.A1(_11251_),
    .A2(_11261_),
    .B1(_11253_),
    .C1(_11262_),
    .D1(_11149_),
    .Y(_11263_));
 sky130_fd_sc_hd__nand3_4 _33823_ (.A(_11258_),
    .B(_11260_),
    .C(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__a21o_4 _33824_ (.A1(_11149_),
    .A2(_11262_),
    .B1(_11257_),
    .X(_11265_));
 sky130_fd_sc_hd__a31oi_4 _33825_ (.A1(_10758_),
    .A2(_10868_),
    .A3(_10859_),
    .B1(_10878_),
    .Y(_11266_));
 sky130_fd_sc_hd__nand3_4 _33826_ (.A(_11257_),
    .B(_11149_),
    .C(_11262_),
    .Y(_11267_));
 sky130_fd_sc_hd__nand3_4 _33827_ (.A(_11265_),
    .B(_11266_),
    .C(_11267_),
    .Y(_11268_));
 sky130_fd_sc_hd__and2b_1 _33828_ (.A_N(_10808_),
    .B(_10800_),
    .X(_11269_));
 sky130_vsdinv _33829_ (.A(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__a21o_1 _33830_ (.A1(_10875_),
    .A2(_10854_),
    .B1(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__nand3_4 _33831_ (.A(_10875_),
    .B(_10854_),
    .C(_11270_),
    .Y(_11272_));
 sky130_fd_sc_hd__nand2_1 _33832_ (.A(_11271_),
    .B(_11272_),
    .Y(_11273_));
 sky130_fd_sc_hd__and2_1 _33833_ (.A(_11273_),
    .B(_18696_),
    .X(_11274_));
 sky130_fd_sc_hd__buf_4 _33834_ (.A(_10968_),
    .X(_11275_));
 sky130_fd_sc_hd__clkbuf_4 _33835_ (.A(_11275_),
    .X(_11276_));
 sky130_fd_sc_hd__nand3_4 _33836_ (.A(_11271_),
    .B(_11276_),
    .C(_11272_),
    .Y(_11277_));
 sky130_vsdinv _33837_ (.A(_11277_),
    .Y(_11278_));
 sky130_fd_sc_hd__o2bb2ai_2 _33838_ (.A1_N(_11264_),
    .A2_N(_11268_),
    .B1(_11274_),
    .B2(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__a21boi_2 _33839_ (.A1(_10884_),
    .A2(_10896_),
    .B1_N(_10872_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand2_1 _33840_ (.A(_11273_),
    .B(_11276_),
    .Y(_11281_));
 sky130_fd_sc_hd__nand3_1 _33841_ (.A(_11271_),
    .B(_18696_),
    .C(_11272_),
    .Y(_11282_));
 sky130_fd_sc_hd__nand2_1 _33842_ (.A(_11281_),
    .B(_11282_),
    .Y(_11283_));
 sky130_fd_sc_hd__nand3_2 _33843_ (.A(_11283_),
    .B(_11268_),
    .C(_11264_),
    .Y(_11284_));
 sky130_fd_sc_hd__nand3_4 _33844_ (.A(_11279_),
    .B(_11280_),
    .C(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__nand2_1 _33845_ (.A(_11273_),
    .B(_18696_),
    .Y(_11286_));
 sky130_fd_sc_hd__nand2_4 _33846_ (.A(_11286_),
    .B(_11277_),
    .Y(_11287_));
 sky130_fd_sc_hd__a21o_1 _33847_ (.A1(_11268_),
    .A2(_11264_),
    .B1(_11287_),
    .X(_11288_));
 sky130_fd_sc_hd__nand2_1 _33848_ (.A(_10884_),
    .B(_10896_),
    .Y(_11289_));
 sky130_fd_sc_hd__nand2_1 _33849_ (.A(_11289_),
    .B(_10872_),
    .Y(_11290_));
 sky130_fd_sc_hd__nand3_2 _33850_ (.A(_11287_),
    .B(_11268_),
    .C(_11264_),
    .Y(_11291_));
 sky130_fd_sc_hd__nand3_4 _33851_ (.A(_11288_),
    .B(_11290_),
    .C(_11291_),
    .Y(_11292_));
 sky130_fd_sc_hd__o2bb2ai_2 _33852_ (.A1_N(_11285_),
    .A2_N(_11292_),
    .B1(_10886_),
    .B2(_10888_),
    .Y(_11293_));
 sky130_fd_sc_hd__nand3_4 _33853_ (.A(_11292_),
    .B(_10895_),
    .C(_11285_),
    .Y(_11294_));
 sky130_fd_sc_hd__nand2_1 _33854_ (.A(_10898_),
    .B(_10534_),
    .Y(_11295_));
 sky130_fd_sc_hd__nand2_2 _33855_ (.A(_11295_),
    .B(_10904_),
    .Y(_11296_));
 sky130_fd_sc_hd__a21o_2 _33856_ (.A1(_11293_),
    .A2(_11294_),
    .B1(_11296_),
    .X(_11297_));
 sky130_fd_sc_hd__nand3_4 _33857_ (.A(_11293_),
    .B(_11294_),
    .C(_11296_),
    .Y(_11298_));
 sky130_fd_sc_hd__nand2_4 _33858_ (.A(_11297_),
    .B(_11298_),
    .Y(_11299_));
 sky130_fd_sc_hd__o2111ai_4 _33859_ (.A1(_10906_),
    .A2(_10911_),
    .B1(_10548_),
    .C1(_10544_),
    .D1(_10912_),
    .Y(_11300_));
 sky130_fd_sc_hd__nor3_4 _33860_ (.A(_10200_),
    .B(_11300_),
    .C(_09872_),
    .Y(_11301_));
 sky130_fd_sc_hd__o2111ai_4 _33861_ (.A1(_06597_),
    .A2(_06416_),
    .B1(_08677_),
    .C1(_06600_),
    .D1(_11301_),
    .Y(_11302_));
 sky130_fd_sc_hd__nor2_2 _33862_ (.A(_10200_),
    .B(_11300_),
    .Y(_11303_));
 sky130_vsdinv _33863_ (.A(_10548_),
    .Y(_11304_));
 sky130_fd_sc_hd__a2bb2oi_4 _33864_ (.A1_N(_10906_),
    .A2_N(_10911_),
    .B1(_10912_),
    .B2(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__o21ai_4 _33865_ (.A1(_10204_),
    .A2(_11300_),
    .B1(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__a21oi_4 _33866_ (.A1(_09875_),
    .A2(_11303_),
    .B1(_11306_),
    .Y(_11307_));
 sky130_fd_sc_hd__nand2_1 _33867_ (.A(_08681_),
    .B(_11301_),
    .Y(_11308_));
 sky130_fd_sc_hd__nand3_4 _33868_ (.A(_11302_),
    .B(_11307_),
    .C(_11308_),
    .Y(_11309_));
 sky130_fd_sc_hd__xnor2_2 _33869_ (.A(_11299_),
    .B(_11309_),
    .Y(_02651_));
 sky130_vsdinv _33870_ (.A(_11194_),
    .Y(_11310_));
 sky130_fd_sc_hd__nor2_8 _33871_ (.A(_11310_),
    .B(_11202_),
    .Y(_11311_));
 sky130_fd_sc_hd__nand2_2 _33872_ (.A(_11261_),
    .B(_11255_),
    .Y(_11312_));
 sky130_fd_sc_hd__nor2_4 _33873_ (.A(_11311_),
    .B(_11312_),
    .Y(_11313_));
 sky130_vsdinv _33874_ (.A(_11311_),
    .Y(_11314_));
 sky130_fd_sc_hd__and2_4 _33875_ (.A(_11261_),
    .B(_11255_),
    .X(_11315_));
 sky130_fd_sc_hd__nor2_4 _33876_ (.A(_11314_),
    .B(_11315_),
    .Y(_11316_));
 sky130_fd_sc_hd__o21ai_2 _33877_ (.A1(_11147_),
    .A2(_11052_),
    .B1(_11143_),
    .Y(_11317_));
 sky130_fd_sc_hd__o21ai_2 _33878_ (.A1(_11045_),
    .A2(_10958_),
    .B1(_10955_),
    .Y(_11318_));
 sky130_fd_sc_hd__o21ai_4 _33879_ (.A1(_10958_),
    .A2(_10959_),
    .B1(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__o21ai_4 _33880_ (.A1(_11032_),
    .A2(_11319_),
    .B1(_11049_),
    .Y(_11320_));
 sky130_fd_sc_hd__nand3_4 _33881_ (.A(_10961_),
    .B(_10962_),
    .C(_20170_),
    .Y(_11321_));
 sky130_fd_sc_hd__nor2_2 _33882_ (.A(_07901_),
    .B(_11321_),
    .Y(_11322_));
 sky130_fd_sc_hd__a22oi_4 _33883_ (.A1(_10972_),
    .A2(_20171_),
    .B1(_05132_),
    .B2(_10973_),
    .Y(_11323_));
 sky130_fd_sc_hd__nand2_4 _33884_ (.A(_10577_),
    .B(_05451_),
    .Y(_11324_));
 sky130_fd_sc_hd__o21ai_2 _33885_ (.A1(_11322_),
    .A2(_11323_),
    .B1(_11324_),
    .Y(_11325_));
 sky130_vsdinv _33886_ (.A(_11324_),
    .Y(_11326_));
 sky130_fd_sc_hd__o2bb2ai_4 _33887_ (.A1_N(_19829_),
    .A2_N(_05179_),
    .B1(_07901_),
    .B2(_10967_),
    .Y(_11327_));
 sky130_fd_sc_hd__o211ai_4 _33888_ (.A1(_20175_),
    .A2(_11321_),
    .B1(_11326_),
    .C1(_11327_),
    .Y(_11328_));
 sky130_fd_sc_hd__o22ai_4 _33889_ (.A1(_20178_),
    .A2(_10963_),
    .B1(_10965_),
    .B2(_10974_),
    .Y(_11329_));
 sky130_fd_sc_hd__nand3_4 _33890_ (.A(_11325_),
    .B(_11328_),
    .C(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__o21ai_2 _33891_ (.A1(_11322_),
    .A2(_11323_),
    .B1(_11326_),
    .Y(_11331_));
 sky130_fd_sc_hd__nand3b_2 _33892_ (.A_N(_11322_),
    .B(_11324_),
    .C(_11327_),
    .Y(_11332_));
 sky130_fd_sc_hd__o21ai_1 _33893_ (.A1(_05415_),
    .A2(_10963_),
    .B1(_10965_),
    .Y(_11333_));
 sky130_fd_sc_hd__nand2_2 _33894_ (.A(_11333_),
    .B(_10969_),
    .Y(_11334_));
 sky130_fd_sc_hd__nand3_4 _33895_ (.A(_11331_),
    .B(_11332_),
    .C(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__buf_2 _33896_ (.A(_10983_),
    .X(_11336_));
 sky130_fd_sc_hd__nand2_2 _33897_ (.A(_19835_),
    .B(_05283_),
    .Y(_11337_));
 sky130_fd_sc_hd__nand2_2 _33898_ (.A(_10000_),
    .B(_05388_),
    .Y(_11338_));
 sky130_fd_sc_hd__nand2_2 _33899_ (.A(_11337_),
    .B(_11338_),
    .Y(_11339_));
 sky130_fd_sc_hd__o21ai_1 _33900_ (.A1(_07752_),
    .A2(_11336_),
    .B1(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__nand2_4 _33901_ (.A(_19843_),
    .B(_05684_),
    .Y(_11341_));
 sky130_vsdinv _33902_ (.A(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__nand2_1 _33903_ (.A(_11340_),
    .B(_11342_),
    .Y(_11343_));
 sky130_vsdinv _33904_ (.A(_11343_),
    .Y(_11344_));
 sky130_fd_sc_hd__nor2_2 _33905_ (.A(_07752_),
    .B(_10987_),
    .Y(_11345_));
 sky130_fd_sc_hd__nand3b_2 _33906_ (.A_N(_11345_),
    .B(_11339_),
    .C(_11341_),
    .Y(_11346_));
 sky130_vsdinv _33907_ (.A(_11346_),
    .Y(_11347_));
 sky130_fd_sc_hd__o2bb2ai_2 _33908_ (.A1_N(_11330_),
    .A2_N(_11335_),
    .B1(_11344_),
    .B2(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__nor2_1 _33909_ (.A(_10965_),
    .B(_10964_),
    .Y(_11349_));
 sky130_fd_sc_hd__a21oi_2 _33910_ (.A1(_11349_),
    .A2(_10969_),
    .B1(_10976_),
    .Y(_11350_));
 sky130_fd_sc_hd__a21oi_2 _33911_ (.A1(_10978_),
    .A2(_10996_),
    .B1(_11350_),
    .Y(_11351_));
 sky130_fd_sc_hd__nand2_2 _33912_ (.A(_11346_),
    .B(_11343_),
    .Y(_11352_));
 sky130_fd_sc_hd__nand3b_2 _33913_ (.A_N(_11352_),
    .B(_11335_),
    .C(_11330_),
    .Y(_11353_));
 sky130_fd_sc_hd__nand3_4 _33914_ (.A(_11348_),
    .B(_11351_),
    .C(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__a21o_1 _33915_ (.A1(_10978_),
    .A2(_10996_),
    .B1(_11350_),
    .X(_11355_));
 sky130_fd_sc_hd__a21oi_4 _33916_ (.A1(_11337_),
    .A2(_11338_),
    .B1(_11341_),
    .Y(_11356_));
 sky130_fd_sc_hd__o21a_1 _33917_ (.A1(_11337_),
    .A2(_11338_),
    .B1(_11356_),
    .X(_11357_));
 sky130_vsdinv _33918_ (.A(_11340_),
    .Y(_11358_));
 sky130_fd_sc_hd__nor2_1 _33919_ (.A(_11342_),
    .B(_11358_),
    .Y(_11359_));
 sky130_fd_sc_hd__o2bb2ai_1 _33920_ (.A1_N(_11330_),
    .A2_N(_11335_),
    .B1(_11357_),
    .B2(_11359_),
    .Y(_11360_));
 sky130_fd_sc_hd__nand3_2 _33921_ (.A(_11335_),
    .B(_11330_),
    .C(_11352_),
    .Y(_11361_));
 sky130_fd_sc_hd__nand3_4 _33922_ (.A(_11355_),
    .B(_11360_),
    .C(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__buf_4 _33923_ (.A(_08800_),
    .X(_11363_));
 sky130_fd_sc_hd__nand2_2 _33924_ (.A(_11008_),
    .B(_05799_),
    .Y(_11364_));
 sky130_fd_sc_hd__a21o_1 _33925_ (.A1(_11363_),
    .A2(_20153_),
    .B1(_11364_),
    .X(_11365_));
 sky130_fd_sc_hd__clkbuf_4 _33926_ (.A(_11008_),
    .X(_11366_));
 sky130_fd_sc_hd__nand2_2 _33927_ (.A(_10553_),
    .B(_05991_),
    .Y(_11367_));
 sky130_fd_sc_hd__a21o_1 _33928_ (.A1(_11366_),
    .A2(_20157_),
    .B1(_11367_),
    .X(_11368_));
 sky130_fd_sc_hd__nand2_2 _33929_ (.A(_08802_),
    .B(_10611_),
    .Y(_11369_));
 sky130_fd_sc_hd__nand3_4 _33930_ (.A(_11365_),
    .B(_11368_),
    .C(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__buf_6 _33931_ (.A(_19850_),
    .X(_11371_));
 sky130_fd_sc_hd__nand3b_4 _33932_ (.A_N(_11364_),
    .B(_11371_),
    .C(_05832_),
    .Y(_11372_));
 sky130_vsdinv _33933_ (.A(_11369_),
    .Y(_11373_));
 sky130_fd_sc_hd__nand2_4 _33934_ (.A(_11364_),
    .B(_11367_),
    .Y(_11374_));
 sky130_fd_sc_hd__nand3_4 _33935_ (.A(_11372_),
    .B(_11373_),
    .C(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__nor2_1 _33936_ (.A(_10980_),
    .B(_10984_),
    .Y(_11376_));
 sky130_fd_sc_hd__o2bb2ai_2 _33937_ (.A1_N(_11370_),
    .A2_N(_11375_),
    .B1(_10981_),
    .B2(_11376_),
    .Y(_11377_));
 sky130_fd_sc_hd__o22ai_4 _33938_ (.A1(_05863_),
    .A2(_11336_),
    .B1(_10979_),
    .B2(_10981_),
    .Y(_11378_));
 sky130_fd_sc_hd__nand3_4 _33939_ (.A(_11370_),
    .B(_11375_),
    .C(_11378_),
    .Y(_11379_));
 sky130_fd_sc_hd__o21a_2 _33940_ (.A1(_11009_),
    .A2(_11006_),
    .B1(_11016_),
    .X(_11380_));
 sky130_vsdinv _33941_ (.A(_11380_),
    .Y(_11381_));
 sky130_fd_sc_hd__a21oi_4 _33942_ (.A1(_11377_),
    .A2(_11379_),
    .B1(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__and3_1 _33943_ (.A(_11381_),
    .B(_11377_),
    .C(_11379_),
    .X(_11383_));
 sky130_fd_sc_hd__o2bb2ai_2 _33944_ (.A1_N(_11354_),
    .A2_N(_11362_),
    .B1(_11382_),
    .B2(_11383_),
    .Y(_11384_));
 sky130_fd_sc_hd__o2bb2ai_2 _33945_ (.A1_N(_11028_),
    .A2_N(_11004_),
    .B1(_11033_),
    .B2(_11037_),
    .Y(_11385_));
 sky130_fd_sc_hd__a21oi_4 _33946_ (.A1(_11370_),
    .A2(_11375_),
    .B1(_11378_),
    .Y(_11386_));
 sky130_fd_sc_hd__nor2_4 _33947_ (.A(_11380_),
    .B(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__a21oi_4 _33948_ (.A1(_11379_),
    .A2(_11387_),
    .B1(_11382_),
    .Y(_11388_));
 sky130_fd_sc_hd__nand3_4 _33949_ (.A(_11388_),
    .B(_11354_),
    .C(_11362_),
    .Y(_11389_));
 sky130_fd_sc_hd__nand3_4 _33950_ (.A(_11384_),
    .B(_11385_),
    .C(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__nand2_1 _33951_ (.A(_11362_),
    .B(_11354_),
    .Y(_11391_));
 sky130_fd_sc_hd__nand2_1 _33952_ (.A(_11391_),
    .B(_11388_),
    .Y(_11392_));
 sky130_fd_sc_hd__a21boi_4 _33953_ (.A1(_11028_),
    .A2(_11004_),
    .B1_N(_10998_),
    .Y(_11393_));
 sky130_fd_sc_hd__o211ai_2 _33954_ (.A1(_11382_),
    .A2(_11383_),
    .B1(_11354_),
    .C1(_11362_),
    .Y(_11394_));
 sky130_fd_sc_hd__nand3_4 _33955_ (.A(_11392_),
    .B(_11393_),
    .C(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__buf_6 _33956_ (.A(_10610_),
    .X(_11396_));
 sky130_fd_sc_hd__a22oi_4 _33957_ (.A1(_11396_),
    .A2(_20147_),
    .B1(_10918_),
    .B2(_20143_),
    .Y(_11397_));
 sky130_fd_sc_hd__nand3_4 _33958_ (.A(_10610_),
    .B(_10620_),
    .C(_05823_),
    .Y(_11398_));
 sky130_fd_sc_hd__nor2_4 _33959_ (.A(_05813_),
    .B(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_4 _33960_ (.A(_07967_),
    .B(_07185_),
    .Y(_11400_));
 sky130_vsdinv _33961_ (.A(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__o21ai_2 _33962_ (.A1(_11397_),
    .A2(_11399_),
    .B1(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__a21oi_4 _33963_ (.A1(_10927_),
    .A2(_10923_),
    .B1(_10921_),
    .Y(_11403_));
 sky130_fd_sc_hd__a22o_1 _33964_ (.A1(_10917_),
    .A2(_10919_),
    .B1(_10926_),
    .B2(_08008_),
    .X(_11404_));
 sky130_fd_sc_hd__o211ai_2 _33965_ (.A1(_06308_),
    .A2(_11398_),
    .B1(_11400_),
    .C1(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__nand3_4 _33966_ (.A(_11402_),
    .B(_11403_),
    .C(_11405_),
    .Y(_11406_));
 sky130_fd_sc_hd__o21ai_2 _33967_ (.A1(_11397_),
    .A2(_11399_),
    .B1(_11400_),
    .Y(_11407_));
 sky130_fd_sc_hd__o22ai_4 _33968_ (.A1(_06298_),
    .A2(_10619_),
    .B1(_10922_),
    .B2(_10920_),
    .Y(_11408_));
 sky130_fd_sc_hd__o211ai_2 _33969_ (.A1(_06308_),
    .A2(_11398_),
    .B1(_11401_),
    .C1(_11404_),
    .Y(_11409_));
 sky130_fd_sc_hd__nand3_4 _33970_ (.A(_11407_),
    .B(_11408_),
    .C(_11409_),
    .Y(_11410_));
 sky130_fd_sc_hd__nand2_2 _33971_ (.A(_10934_),
    .B(_06143_),
    .Y(_11411_));
 sky130_fd_sc_hd__nand2_2 _33972_ (.A(_10944_),
    .B(_07003_),
    .Y(_11412_));
 sky130_fd_sc_hd__nor2_1 _33973_ (.A(_11411_),
    .B(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__nand2_4 _33974_ (.A(_19877_),
    .B(_20130_),
    .Y(_11414_));
 sky130_fd_sc_hd__nand2_1 _33975_ (.A(_11411_),
    .B(_11412_),
    .Y(_11415_));
 sky130_fd_sc_hd__nand3b_2 _33976_ (.A_N(_11413_),
    .B(_11414_),
    .C(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__a22oi_4 _33977_ (.A1(_10935_),
    .A2(_20136_),
    .B1(_10936_),
    .B2(_20134_),
    .Y(_11417_));
 sky130_fd_sc_hd__buf_2 _33978_ (.A(_11413_),
    .X(_11418_));
 sky130_vsdinv _33979_ (.A(_11414_),
    .Y(_11419_));
 sky130_fd_sc_hd__o21ai_1 _33980_ (.A1(_11417_),
    .A2(_11418_),
    .B1(_11419_),
    .Y(_11420_));
 sky130_fd_sc_hd__nand2_2 _33981_ (.A(_11416_),
    .B(_11420_),
    .Y(_11421_));
 sky130_fd_sc_hd__a21oi_2 _33982_ (.A1(_11406_),
    .A2(_11410_),
    .B1(_11421_),
    .Y(_11422_));
 sky130_fd_sc_hd__nor3_1 _33983_ (.A(_11419_),
    .B(_11417_),
    .C(_11418_),
    .Y(_11423_));
 sky130_fd_sc_hd__o21a_1 _33984_ (.A1(_11417_),
    .A2(_11418_),
    .B1(_11419_),
    .X(_11424_));
 sky130_fd_sc_hd__o211a_1 _33985_ (.A1(_11423_),
    .A2(_11424_),
    .B1(_11410_),
    .C1(_11406_),
    .X(_11425_));
 sky130_fd_sc_hd__o21ai_4 _33986_ (.A1(_11023_),
    .A2(_11024_),
    .B1(_11021_),
    .Y(_11426_));
 sky130_fd_sc_hd__o21bai_4 _33987_ (.A1(_11422_),
    .A2(_11425_),
    .B1_N(_11426_),
    .Y(_11427_));
 sky130_fd_sc_hd__o21a_1 _33988_ (.A1(_11417_),
    .A2(_11418_),
    .B1(_11414_),
    .X(_11428_));
 sky130_fd_sc_hd__nor3_4 _33989_ (.A(_11414_),
    .B(_11417_),
    .C(_11418_),
    .Y(_11429_));
 sky130_fd_sc_hd__o2bb2ai_4 _33990_ (.A1_N(_11410_),
    .A2_N(_11406_),
    .B1(_11428_),
    .B2(_11429_),
    .Y(_11430_));
 sky130_fd_sc_hd__nand3_4 _33991_ (.A(_11406_),
    .B(_11421_),
    .C(_11410_),
    .Y(_11431_));
 sky130_fd_sc_hd__nand3_4 _33992_ (.A(_11430_),
    .B(_11426_),
    .C(_11431_),
    .Y(_11432_));
 sky130_fd_sc_hd__nand2_1 _33993_ (.A(_10929_),
    .B(_10949_),
    .Y(_11433_));
 sky130_fd_sc_hd__nand2_4 _33994_ (.A(_11433_),
    .B(_10933_),
    .Y(_11434_));
 sky130_fd_sc_hd__nand3_2 _33995_ (.A(_11427_),
    .B(_11432_),
    .C(_11434_),
    .Y(_11435_));
 sky130_vsdinv _33996_ (.A(_11435_),
    .Y(_11436_));
 sky130_fd_sc_hd__a21oi_4 _33997_ (.A1(_11427_),
    .A2(_11432_),
    .B1(_11434_),
    .Y(_11437_));
 sky130_fd_sc_hd__o2bb2ai_2 _33998_ (.A1_N(_11390_),
    .A2_N(_11395_),
    .B1(_11436_),
    .B2(_11437_),
    .Y(_11438_));
 sky130_vsdinv _33999_ (.A(_11434_),
    .Y(_11439_));
 sky130_fd_sc_hd__a21oi_4 _34000_ (.A1(_11430_),
    .A2(_11431_),
    .B1(_11426_),
    .Y(_11440_));
 sky130_fd_sc_hd__nor2_2 _34001_ (.A(_11439_),
    .B(_11440_),
    .Y(_11441_));
 sky130_fd_sc_hd__a21oi_4 _34002_ (.A1(_11432_),
    .A2(_11441_),
    .B1(_11437_),
    .Y(_11442_));
 sky130_fd_sc_hd__nand3_4 _34003_ (.A(_11442_),
    .B(_11395_),
    .C(_11390_),
    .Y(_11443_));
 sky130_fd_sc_hd__nand3_4 _34004_ (.A(_11320_),
    .B(_11438_),
    .C(_11443_),
    .Y(_11444_));
 sky130_fd_sc_hd__a21oi_4 _34005_ (.A1(_11044_),
    .A2(_11048_),
    .B1(_11040_),
    .Y(_11445_));
 sky130_fd_sc_hd__nand2_1 _34006_ (.A(_11395_),
    .B(_11390_),
    .Y(_11446_));
 sky130_fd_sc_hd__nand2_1 _34007_ (.A(_11446_),
    .B(_11442_),
    .Y(_11447_));
 sky130_vsdinv _34008_ (.A(_10929_),
    .Y(_11448_));
 sky130_fd_sc_hd__and3_1 _34009_ (.A(_10933_),
    .B(_10943_),
    .C(_10948_),
    .X(_11449_));
 sky130_fd_sc_hd__and3_1 _34010_ (.A(_11430_),
    .B(_11426_),
    .C(_11431_),
    .X(_11450_));
 sky130_fd_sc_hd__o22ai_2 _34011_ (.A1(_11448_),
    .A2(_11449_),
    .B1(_11440_),
    .B2(_11450_),
    .Y(_11451_));
 sky130_fd_sc_hd__nand2_2 _34012_ (.A(_11451_),
    .B(_11435_),
    .Y(_11452_));
 sky130_fd_sc_hd__nand3_2 _34013_ (.A(_11395_),
    .B(_11452_),
    .C(_11390_),
    .Y(_11453_));
 sky130_fd_sc_hd__nand3_4 _34014_ (.A(_11445_),
    .B(_11447_),
    .C(_11453_),
    .Y(_11454_));
 sky130_fd_sc_hd__buf_4 _34015_ (.A(_07295_),
    .X(_11455_));
 sky130_fd_sc_hd__a22oi_4 _34016_ (.A1(_19882_),
    .A2(_20127_),
    .B1(_11455_),
    .B2(_07568_),
    .Y(_11456_));
 sky130_fd_sc_hd__buf_6 _34017_ (.A(_08040_),
    .X(_11457_));
 sky130_fd_sc_hd__nand3_4 _34018_ (.A(_11092_),
    .B(_19887_),
    .C(_07258_),
    .Y(_11458_));
 sky130_fd_sc_hd__nor2_4 _34019_ (.A(_11457_),
    .B(_11458_),
    .Y(_11459_));
 sky130_fd_sc_hd__nand2_2 _34020_ (.A(_06641_),
    .B(_07726_),
    .Y(_11460_));
 sky130_fd_sc_hd__o21ai_2 _34021_ (.A1(_11456_),
    .A2(_11459_),
    .B1(_11460_),
    .Y(_11461_));
 sky130_vsdinv _34022_ (.A(_11460_),
    .Y(_11462_));
 sky130_fd_sc_hd__clkbuf_4 _34023_ (.A(_07088_),
    .X(_11463_));
 sky130_fd_sc_hd__a22o_2 _34024_ (.A1(_11463_),
    .A2(_10350_),
    .B1(_11455_),
    .B2(_07568_),
    .X(_11464_));
 sky130_fd_sc_hd__o211ai_4 _34025_ (.A1(_11457_),
    .A2(_11458_),
    .B1(_11462_),
    .C1(_11464_),
    .Y(_11465_));
 sky130_fd_sc_hd__o21ai_2 _34026_ (.A1(_10942_),
    .A2(_10937_),
    .B1(_10946_),
    .Y(_11466_));
 sky130_fd_sc_hd__nand3_4 _34027_ (.A(_11461_),
    .B(_11465_),
    .C(_11466_),
    .Y(_11467_));
 sky130_fd_sc_hd__o21ai_2 _34028_ (.A1(_11456_),
    .A2(_11459_),
    .B1(_11462_),
    .Y(_11468_));
 sky130_fd_sc_hd__o21ai_1 _34029_ (.A1(_10938_),
    .A2(_10939_),
    .B1(_10942_),
    .Y(_11469_));
 sky130_fd_sc_hd__nand2_1 _34030_ (.A(_11469_),
    .B(_10947_),
    .Y(_11470_));
 sky130_fd_sc_hd__o211ai_4 _34031_ (.A1(_11457_),
    .A2(_11458_),
    .B1(_11460_),
    .C1(_11464_),
    .Y(_11471_));
 sky130_fd_sc_hd__nand3_4 _34032_ (.A(_11468_),
    .B(_11470_),
    .C(_11471_),
    .Y(_11472_));
 sky130_fd_sc_hd__nor2_4 _34033_ (.A(_11099_),
    .B(_11097_),
    .Y(_11473_));
 sky130_fd_sc_hd__o2bb2ai_4 _34034_ (.A1_N(_11467_),
    .A2_N(_11472_),
    .B1(_11095_),
    .B2(_11473_),
    .Y(_11474_));
 sky130_fd_sc_hd__nor2_2 _34035_ (.A(_11095_),
    .B(_11473_),
    .Y(_11475_));
 sky130_fd_sc_hd__nand3_4 _34036_ (.A(_11467_),
    .B(_11472_),
    .C(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__nand2_4 _34037_ (.A(_11116_),
    .B(_11111_),
    .Y(_11477_));
 sky130_fd_sc_hd__a21oi_4 _34038_ (.A1(_11474_),
    .A2(_11476_),
    .B1(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__a21oi_2 _34039_ (.A1(_10669_),
    .A2(_10672_),
    .B1(_10678_),
    .Y(_11479_));
 sky130_fd_sc_hd__a31oi_2 _34040_ (.A1(_11100_),
    .A2(_11102_),
    .A3(_11105_),
    .B1(_11479_),
    .Y(_11480_));
 sky130_vsdinv _34041_ (.A(_11111_),
    .Y(_11481_));
 sky130_fd_sc_hd__o211a_4 _34042_ (.A1(_11480_),
    .A2(_11481_),
    .B1(_11476_),
    .C1(_11474_),
    .X(_11482_));
 sky130_fd_sc_hd__a21o_1 _34043_ (.A1(_11063_),
    .A2(_11065_),
    .B1(_11060_),
    .X(_11483_));
 sky130_fd_sc_hd__nand3_4 _34044_ (.A(_19893_),
    .B(_06359_),
    .C(_20114_),
    .Y(_11484_));
 sky130_fd_sc_hd__nor2_8 _34045_ (.A(_10340_),
    .B(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__clkbuf_4 _34046_ (.A(_07922_),
    .X(_11486_));
 sky130_fd_sc_hd__buf_4 _34047_ (.A(_07722_),
    .X(_11487_));
 sky130_fd_sc_hd__a22o_2 _34048_ (.A1(_11486_),
    .A2(_07561_),
    .B1(_07115_),
    .B2(_11487_),
    .X(_11488_));
 sky130_fd_sc_hd__nand2_2 _34049_ (.A(net505),
    .B(_20107_),
    .Y(_11489_));
 sky130_vsdinv _34050_ (.A(_11489_),
    .Y(_11490_));
 sky130_fd_sc_hd__nand3b_2 _34051_ (.A_N(_11485_),
    .B(_11488_),
    .C(_11490_),
    .Y(_11491_));
 sky130_fd_sc_hd__buf_4 _34052_ (.A(_08056_),
    .X(_11492_));
 sky130_fd_sc_hd__a22oi_4 _34053_ (.A1(net444),
    .A2(_09921_),
    .B1(_10351_),
    .B2(_11492_),
    .Y(_11493_));
 sky130_fd_sc_hd__o21ai_2 _34054_ (.A1(_11493_),
    .A2(_11485_),
    .B1(_11489_),
    .Y(_11494_));
 sky130_fd_sc_hd__nand3_4 _34055_ (.A(_11483_),
    .B(_11491_),
    .C(_11494_),
    .Y(_11495_));
 sky130_vsdinv _34056_ (.A(_11495_),
    .Y(_11496_));
 sky130_fd_sc_hd__o21ai_2 _34057_ (.A1(_11493_),
    .A2(_11485_),
    .B1(_11490_),
    .Y(_11497_));
 sky130_fd_sc_hd__a21oi_2 _34058_ (.A1(_11063_),
    .A2(_11065_),
    .B1(_11060_),
    .Y(_11498_));
 sky130_fd_sc_hd__o211ai_2 _34059_ (.A1(_10824_),
    .A2(_11484_),
    .B1(_11489_),
    .C1(_11488_),
    .Y(_11499_));
 sky130_fd_sc_hd__nand3_4 _34060_ (.A(_11497_),
    .B(_11498_),
    .C(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__a22oi_4 _34061_ (.A1(_10337_),
    .A2(_11078_),
    .B1(_10338_),
    .B2(_20102_),
    .Y(_11501_));
 sky130_fd_sc_hd__and4_1 _34062_ (.A(_06048_),
    .B(_06049_),
    .C(_10811_),
    .D(_20105_),
    .X(_11502_));
 sky130_fd_sc_hd__buf_4 _34063_ (.A(_20096_),
    .X(_11503_));
 sky130_fd_sc_hd__nand2_2 _34064_ (.A(_05953_),
    .B(_11503_),
    .Y(_11504_));
 sky130_vsdinv _34065_ (.A(_11504_),
    .Y(_11505_));
 sky130_fd_sc_hd__o21ai_1 _34066_ (.A1(_11501_),
    .A2(_11502_),
    .B1(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__nand2_1 _34067_ (.A(_19906_),
    .B(_10222_),
    .Y(_11507_));
 sky130_fd_sc_hd__nand3b_2 _34068_ (.A_N(_11507_),
    .B(_19903_),
    .C(_11085_),
    .Y(_11508_));
 sky130_fd_sc_hd__a22o_1 _34069_ (.A1(_06119_),
    .A2(_20105_),
    .B1(_10347_),
    .B2(_09044_),
    .X(_11509_));
 sky130_fd_sc_hd__nand3_1 _34070_ (.A(_11508_),
    .B(_11504_),
    .C(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__nand2_1 _34071_ (.A(_11506_),
    .B(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__nand2_2 _34072_ (.A(_11500_),
    .B(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__a21o_1 _34073_ (.A1(_11495_),
    .A2(_11500_),
    .B1(_11511_),
    .X(_11513_));
 sky130_fd_sc_hd__o21ai_4 _34074_ (.A1(_11496_),
    .A2(_11512_),
    .B1(_11513_),
    .Y(_11514_));
 sky130_fd_sc_hd__o21bai_4 _34075_ (.A1(_11478_),
    .A2(_11482_),
    .B1_N(_11514_),
    .Y(_11515_));
 sky130_fd_sc_hd__nand2_1 _34076_ (.A(_10954_),
    .B(_10955_),
    .Y(_11516_));
 sky130_fd_sc_hd__nand2_2 _34077_ (.A(_11516_),
    .B(_10953_),
    .Y(_11517_));
 sky130_fd_sc_hd__a21o_1 _34078_ (.A1(_11476_),
    .A2(_11474_),
    .B1(_11477_),
    .X(_11518_));
 sky130_fd_sc_hd__nand3_4 _34079_ (.A(_11477_),
    .B(_11476_),
    .C(_11474_),
    .Y(_11519_));
 sky130_fd_sc_hd__nand3_4 _34080_ (.A(_11518_),
    .B(_11519_),
    .C(_11514_),
    .Y(_11520_));
 sky130_fd_sc_hd__o21a_2 _34081_ (.A1(_11129_),
    .A2(_11120_),
    .B1(_11125_),
    .X(_11521_));
 sky130_fd_sc_hd__a31oi_4 _34082_ (.A1(_11515_),
    .A2(_11517_),
    .A3(_11520_),
    .B1(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__o21ai_2 _34083_ (.A1(_11478_),
    .A2(_11482_),
    .B1(_11514_),
    .Y(_11523_));
 sky130_fd_sc_hd__o21ai_2 _34084_ (.A1(_10955_),
    .A2(_11045_),
    .B1(_10954_),
    .Y(_11524_));
 sky130_fd_sc_hd__nand3b_2 _34085_ (.A_N(_11514_),
    .B(_11518_),
    .C(_11519_),
    .Y(_11525_));
 sky130_fd_sc_hd__nand3_4 _34086_ (.A(_11523_),
    .B(_11524_),
    .C(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__nand2_1 _34087_ (.A(_11522_),
    .B(_11526_),
    .Y(_11527_));
 sky130_vsdinv _34088_ (.A(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__nand3_4 _34089_ (.A(_11515_),
    .B(_11517_),
    .C(_11520_),
    .Y(_11529_));
 sky130_fd_sc_hd__o21ai_4 _34090_ (.A1(_11129_),
    .A2(_11120_),
    .B1(_11125_),
    .Y(_11530_));
 sky130_fd_sc_hd__a21oi_4 _34091_ (.A1(_11526_),
    .A2(_11529_),
    .B1(_11530_),
    .Y(_11531_));
 sky130_fd_sc_hd__o2bb2ai_2 _34092_ (.A1_N(_11444_),
    .A2_N(_11454_),
    .B1(_11528_),
    .B2(_11531_),
    .Y(_11532_));
 sky130_fd_sc_hd__a21oi_4 _34093_ (.A1(_11526_),
    .A2(_11522_),
    .B1(_11531_),
    .Y(_11533_));
 sky130_fd_sc_hd__nand3_4 _34094_ (.A(_11533_),
    .B(_11454_),
    .C(_11444_),
    .Y(_11534_));
 sky130_fd_sc_hd__nand3_2 _34095_ (.A(_11317_),
    .B(_11532_),
    .C(_11534_),
    .Y(_11535_));
 sky130_fd_sc_hd__buf_6 _34096_ (.A(_11535_),
    .X(_11536_));
 sky130_fd_sc_hd__nand2_1 _34097_ (.A(_11044_),
    .B(_11049_),
    .Y(_11537_));
 sky130_fd_sc_hd__a22oi_4 _34098_ (.A1(_10660_),
    .A2(_10606_),
    .B1(_11537_),
    .B2(_11319_),
    .Y(_11538_));
 sky130_fd_sc_hd__a22oi_4 _34099_ (.A1(_11050_),
    .A2(_11538_),
    .B1(_11142_),
    .B2(_11140_),
    .Y(_11539_));
 sky130_fd_sc_hd__a21o_1 _34100_ (.A1(_11526_),
    .A2(_11529_),
    .B1(_11530_),
    .X(_11540_));
 sky130_fd_sc_hd__nand2_2 _34101_ (.A(_11540_),
    .B(_11527_),
    .Y(_11541_));
 sky130_fd_sc_hd__nand3_2 _34102_ (.A(_11454_),
    .B(_11541_),
    .C(_11444_),
    .Y(_11542_));
 sky130_fd_sc_hd__a21o_1 _34103_ (.A1(_11454_),
    .A2(_11444_),
    .B1(_11541_),
    .X(_11543_));
 sky130_fd_sc_hd__nand3_4 _34104_ (.A(_11539_),
    .B(_11542_),
    .C(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__nand2_2 _34105_ (.A(_11145_),
    .B(_11137_),
    .Y(_11545_));
 sky130_fd_sc_hd__a21oi_4 _34106_ (.A1(_11233_),
    .A2(_11235_),
    .B1(_11231_),
    .Y(_11546_));
 sky130_vsdinv _34107_ (.A(_11229_),
    .Y(_11547_));
 sky130_fd_sc_hd__a22oi_4 _34108_ (.A1(_06096_),
    .A2(_10814_),
    .B1(_06098_),
    .B2(_09902_),
    .Y(_11548_));
 sky130_vsdinv _34109_ (.A(_09037_),
    .Y(_11549_));
 sky130_fd_sc_hd__nand3_4 _34110_ (.A(_19912_),
    .B(_05608_),
    .C(_11210_),
    .Y(_11550_));
 sky130_fd_sc_hd__nor2_8 _34111_ (.A(_11549_),
    .B(_11550_),
    .Y(_11551_));
 sky130_fd_sc_hd__nand2_2 _34112_ (.A(_19918_),
    .B(_20086_),
    .Y(_11552_));
 sky130_vsdinv _34113_ (.A(_11552_),
    .Y(_11553_));
 sky130_fd_sc_hd__o21ai_2 _34114_ (.A1(_11548_),
    .A2(_11551_),
    .B1(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__o21ai_1 _34115_ (.A1(_11080_),
    .A2(_11081_),
    .B1(_11083_),
    .Y(_11555_));
 sky130_fd_sc_hd__nand2_2 _34116_ (.A(_11555_),
    .B(_11087_),
    .Y(_11556_));
 sky130_fd_sc_hd__buf_6 _34117_ (.A(_11549_),
    .X(_11557_));
 sky130_fd_sc_hd__a22o_2 _34118_ (.A1(_10809_),
    .A2(_10814_),
    .B1(_11206_),
    .B2(_20091_),
    .X(_11558_));
 sky130_fd_sc_hd__o211ai_4 _34119_ (.A1(_11557_),
    .A2(_11550_),
    .B1(_11552_),
    .C1(_11558_),
    .Y(_11559_));
 sky130_fd_sc_hd__nand3_4 _34120_ (.A(_11554_),
    .B(_11556_),
    .C(_11559_),
    .Y(_11560_));
 sky130_fd_sc_hd__o21ai_2 _34121_ (.A1(_11548_),
    .A2(_11551_),
    .B1(_11552_),
    .Y(_11561_));
 sky130_fd_sc_hd__o21ai_2 _34122_ (.A1(_11083_),
    .A2(_11079_),
    .B1(_11086_),
    .Y(_11562_));
 sky130_fd_sc_hd__buf_8 _34123_ (.A(_11549_),
    .X(_11563_));
 sky130_fd_sc_hd__o211ai_4 _34124_ (.A1(_11563_),
    .A2(_11550_),
    .B1(_11553_),
    .C1(_11558_),
    .Y(_11564_));
 sky130_fd_sc_hd__nand3_4 _34125_ (.A(_11561_),
    .B(_11562_),
    .C(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__nor2_4 _34126_ (.A(_11213_),
    .B(_11209_),
    .Y(_11566_));
 sky130_fd_sc_hd__o2bb2ai_4 _34127_ (.A1_N(_11560_),
    .A2_N(_11565_),
    .B1(_11207_),
    .B2(_11566_),
    .Y(_11567_));
 sky130_fd_sc_hd__nor2_2 _34128_ (.A(_11207_),
    .B(_11566_),
    .Y(_11568_));
 sky130_fd_sc_hd__nand3_4 _34129_ (.A(_11560_),
    .B(_11565_),
    .C(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__nand2_4 _34130_ (.A(_11127_),
    .B(_11071_),
    .Y(_11570_));
 sky130_fd_sc_hd__a21oi_4 _34131_ (.A1(_11567_),
    .A2(_11569_),
    .B1(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__and3_1 _34132_ (.A(_11561_),
    .B(_11562_),
    .C(_11564_),
    .X(_11572_));
 sky130_fd_sc_hd__nand2_1 _34133_ (.A(_11560_),
    .B(_11568_),
    .Y(_11573_));
 sky130_fd_sc_hd__o211a_2 _34134_ (.A1(_11572_),
    .A2(_11573_),
    .B1(_11567_),
    .C1(_11570_),
    .X(_11574_));
 sky130_fd_sc_hd__o22ai_4 _34135_ (.A1(_11230_),
    .A2(_11547_),
    .B1(_11571_),
    .B2(_11574_),
    .Y(_11575_));
 sky130_fd_sc_hd__a21o_1 _34136_ (.A1(_11567_),
    .A2(_11569_),
    .B1(_11570_),
    .X(_11576_));
 sky130_fd_sc_hd__nand3_4 _34137_ (.A(_11570_),
    .B(_11567_),
    .C(_11569_),
    .Y(_11577_));
 sky130_fd_sc_hd__nand2_2 _34138_ (.A(_11229_),
    .B(_11217_),
    .Y(_11578_));
 sky130_vsdinv _34139_ (.A(_11578_),
    .Y(_11579_));
 sky130_fd_sc_hd__nand3_2 _34140_ (.A(_11576_),
    .B(_11577_),
    .C(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__nand3_4 _34141_ (.A(_11546_),
    .B(_11575_),
    .C(_11580_),
    .Y(_11581_));
 sky130_fd_sc_hd__o21bai_2 _34142_ (.A1(_11571_),
    .A2(_11574_),
    .B1_N(_11578_),
    .Y(_11582_));
 sky130_vsdinv _34143_ (.A(_11235_),
    .Y(_11583_));
 sky130_fd_sc_hd__o21ai_2 _34144_ (.A1(_11583_),
    .A2(_11228_),
    .B1(_11234_),
    .Y(_11584_));
 sky130_fd_sc_hd__nand3_2 _34145_ (.A(_11576_),
    .B(_11578_),
    .C(_11577_),
    .Y(_11585_));
 sky130_fd_sc_hd__nand3_4 _34146_ (.A(_11582_),
    .B(_11584_),
    .C(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__buf_6 _34147_ (.A(\pcpi_mul.rs1[29] ),
    .X(_11587_));
 sky130_fd_sc_hd__a22oi_4 _34148_ (.A1(_05229_),
    .A2(_09896_),
    .B1(net447),
    .B2(_11587_),
    .Y(_11588_));
 sky130_fd_sc_hd__nor2_4 _34149_ (.A(_11160_),
    .B(_11588_),
    .Y(_11589_));
 sky130_fd_sc_hd__nand2_4 _34150_ (.A(_05229_),
    .B(_20082_),
    .Y(_11590_));
 sky130_fd_sc_hd__nand2_4 _34151_ (.A(net447),
    .B(_20078_),
    .Y(_11591_));
 sky130_fd_sc_hd__or2_1 _34152_ (.A(_11590_),
    .B(_11591_),
    .X(_11592_));
 sky130_fd_sc_hd__nand2_1 _34153_ (.A(_11589_),
    .B(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__a21o_1 _34154_ (.A1(_11162_),
    .A2(_11163_),
    .B1(_11159_),
    .X(_11594_));
 sky130_fd_sc_hd__nor2_8 _34155_ (.A(_11590_),
    .B(_11591_),
    .Y(_11595_));
 sky130_fd_sc_hd__o21ai_2 _34156_ (.A1(_11588_),
    .A2(_11595_),
    .B1(_11168_),
    .Y(_11596_));
 sky130_fd_sc_hd__nand3_4 _34157_ (.A(_11593_),
    .B(_11594_),
    .C(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__nand2_1 _34158_ (.A(_11590_),
    .B(_11591_),
    .Y(_11598_));
 sky130_fd_sc_hd__nand3_2 _34159_ (.A(_11592_),
    .B(_11168_),
    .C(_11598_),
    .Y(_11599_));
 sky130_fd_sc_hd__a21oi_2 _34160_ (.A1(_11162_),
    .A2(_11163_),
    .B1(_11159_),
    .Y(_11600_));
 sky130_fd_sc_hd__o21ai_2 _34161_ (.A1(_11588_),
    .A2(_11595_),
    .B1(_11162_),
    .Y(_11601_));
 sky130_fd_sc_hd__nand3_4 _34162_ (.A(_11599_),
    .B(_11600_),
    .C(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__buf_6 _34163_ (.A(_18686_),
    .X(_11603_));
 sky130_fd_sc_hd__buf_6 _34164_ (.A(_10777_),
    .X(_11604_));
 sky130_fd_sc_hd__a22oi_4 _34165_ (.A1(_11603_),
    .A2(_19935_),
    .B1(_19932_),
    .B2(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__and4_4 _34166_ (.A(_18686_),
    .B(_05140_),
    .C(_05142_),
    .D(_10778_),
    .X(_11606_));
 sky130_fd_sc_hd__buf_6 _34167_ (.A(_11174_),
    .X(_11607_));
 sky130_fd_sc_hd__nand2_2 _34168_ (.A(_19929_),
    .B(_11607_),
    .Y(_11608_));
 sky130_fd_sc_hd__o21a_1 _34169_ (.A1(_11605_),
    .A2(_11606_),
    .B1(_11608_),
    .X(_11609_));
 sky130_fd_sc_hd__nor3_4 _34170_ (.A(_11608_),
    .B(_11605_),
    .C(_11606_),
    .Y(_11610_));
 sky130_fd_sc_hd__o2bb2ai_4 _34171_ (.A1_N(_11597_),
    .A2_N(_11602_),
    .B1(_11609_),
    .B2(_11610_),
    .Y(_11611_));
 sky130_fd_sc_hd__nor2_2 _34172_ (.A(_11610_),
    .B(_11609_),
    .Y(_11612_));
 sky130_fd_sc_hd__nand3_4 _34173_ (.A(_11612_),
    .B(_11597_),
    .C(_11602_),
    .Y(_11613_));
 sky130_fd_sc_hd__o21ai_4 _34174_ (.A1(_11186_),
    .A2(_11171_),
    .B1(_11192_),
    .Y(_11614_));
 sky130_fd_sc_hd__a21o_1 _34175_ (.A1(_11611_),
    .A2(_11613_),
    .B1(_11614_),
    .X(_11615_));
 sky130_fd_sc_hd__nand3_4 _34176_ (.A(_11614_),
    .B(_11611_),
    .C(_11613_),
    .Y(_11616_));
 sky130_fd_sc_hd__a21o_2 _34177_ (.A1(_11184_),
    .A2(_11182_),
    .B1(_11175_),
    .X(_11617_));
 sky130_fd_sc_hd__a21oi_4 _34178_ (.A1(_11615_),
    .A2(_11616_),
    .B1(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__a21oi_4 _34179_ (.A1(_11611_),
    .A2(_11613_),
    .B1(_11614_),
    .Y(_11619_));
 sky130_fd_sc_hd__nand2_4 _34180_ (.A(_11616_),
    .B(_11617_),
    .Y(_11620_));
 sky130_fd_sc_hd__nor2_8 _34181_ (.A(_11619_),
    .B(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__o2bb2ai_2 _34182_ (.A1_N(_11581_),
    .A2_N(_11586_),
    .B1(_11618_),
    .B2(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__nor2_4 _34183_ (.A(_11621_),
    .B(_11618_),
    .Y(_11623_));
 sky130_fd_sc_hd__nand3_4 _34184_ (.A(_11623_),
    .B(_11581_),
    .C(_11586_),
    .Y(_11624_));
 sky130_fd_sc_hd__nand3_4 _34185_ (.A(_11545_),
    .B(_11622_),
    .C(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__nand2_1 _34186_ (.A(_11581_),
    .B(_11586_),
    .Y(_11626_));
 sky130_fd_sc_hd__nand2_2 _34187_ (.A(_11626_),
    .B(_11623_),
    .Y(_11627_));
 sky130_fd_sc_hd__a21oi_4 _34188_ (.A1(_11131_),
    .A2(_11138_),
    .B1(_11144_),
    .Y(_11628_));
 sky130_fd_sc_hd__a21o_1 _34189_ (.A1(_11615_),
    .A2(_11616_),
    .B1(_11617_),
    .X(_11629_));
 sky130_fd_sc_hd__o21ai_4 _34190_ (.A1(_11619_),
    .A2(_11620_),
    .B1(_11629_),
    .Y(_11630_));
 sky130_fd_sc_hd__nand3_4 _34191_ (.A(_11630_),
    .B(_11581_),
    .C(_11586_),
    .Y(_11631_));
 sky130_fd_sc_hd__nand3_4 _34192_ (.A(_11627_),
    .B(_11628_),
    .C(_11631_),
    .Y(_11632_));
 sky130_fd_sc_hd__a21oi_4 _34193_ (.A1(_11242_),
    .A2(_11243_),
    .B1(_11240_),
    .Y(_11633_));
 sky130_vsdinv _34194_ (.A(_11633_),
    .Y(_11634_));
 sky130_fd_sc_hd__a21oi_4 _34195_ (.A1(_11625_),
    .A2(_11632_),
    .B1(_11634_),
    .Y(_11635_));
 sky130_fd_sc_hd__buf_2 _34196_ (.A(_11625_),
    .X(_11636_));
 sky130_fd_sc_hd__nand3_4 _34197_ (.A(_11634_),
    .B(_11632_),
    .C(_11636_),
    .Y(_11637_));
 sky130_vsdinv _34198_ (.A(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__o2bb2ai_4 _34199_ (.A1_N(_11536_),
    .A2_N(_11544_),
    .B1(_11635_),
    .B2(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__a31oi_4 _34200_ (.A1(_11627_),
    .A2(_11628_),
    .A3(_11631_),
    .B1(_11633_),
    .Y(_11640_));
 sky130_fd_sc_hd__a21oi_4 _34201_ (.A1(_11636_),
    .A2(_11640_),
    .B1(_11635_),
    .Y(_11641_));
 sky130_fd_sc_hd__nand3_4 _34202_ (.A(_11544_),
    .B(_11641_),
    .C(_11536_),
    .Y(_11642_));
 sky130_fd_sc_hd__a21oi_4 _34203_ (.A1(_11151_),
    .A2(_11153_),
    .B1(_11152_),
    .Y(_11643_));
 sky130_fd_sc_hd__o21ai_4 _34204_ (.A1(_11257_),
    .A2(_11643_),
    .B1(_11262_),
    .Y(_11644_));
 sky130_fd_sc_hd__a21oi_4 _34205_ (.A1(_11639_),
    .A2(_11642_),
    .B1(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__nand2_1 _34206_ (.A(_11532_),
    .B(_11534_),
    .Y(_11646_));
 sky130_fd_sc_hd__nand2_1 _34207_ (.A(_11636_),
    .B(_11632_),
    .Y(_11647_));
 sky130_fd_sc_hd__nand2_1 _34208_ (.A(_11647_),
    .B(_11633_),
    .Y(_11648_));
 sky130_fd_sc_hd__nand2_2 _34209_ (.A(_11648_),
    .B(_11637_),
    .Y(_11649_));
 sky130_fd_sc_hd__a21oi_1 _34210_ (.A1(_11646_),
    .A2(_11539_),
    .B1(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__nand3_1 _34211_ (.A(_11149_),
    .B(_11256_),
    .C(_11253_),
    .Y(_11651_));
 sky130_fd_sc_hd__a21oi_4 _34212_ (.A1(_11544_),
    .A2(_11536_),
    .B1(_11641_),
    .Y(_11652_));
 sky130_fd_sc_hd__a221oi_2 _34213_ (.A1(_11650_),
    .A2(_11536_),
    .B1(_11651_),
    .B2(_11262_),
    .C1(_11652_),
    .Y(_11653_));
 sky130_fd_sc_hd__o22ai_4 _34214_ (.A1(_11313_),
    .A2(_11316_),
    .B1(_11645_),
    .B2(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__a21boi_4 _34215_ (.A1(_11287_),
    .A2(_11268_),
    .B1_N(_11264_),
    .Y(_11655_));
 sky130_fd_sc_hd__and3_1 _34216_ (.A(_11544_),
    .B(_11641_),
    .C(_11535_),
    .X(_11656_));
 sky130_fd_sc_hd__o21a_1 _34217_ (.A1(_11257_),
    .A2(_11643_),
    .B1(_11262_),
    .X(_11657_));
 sky130_fd_sc_hd__o21ai_4 _34218_ (.A1(_11652_),
    .A2(_11656_),
    .B1(_11657_),
    .Y(_11658_));
 sky130_fd_sc_hd__nand3_4 _34219_ (.A(_11644_),
    .B(_11642_),
    .C(_11639_),
    .Y(_11659_));
 sky130_fd_sc_hd__nor2_4 _34220_ (.A(_11313_),
    .B(_11316_),
    .Y(_11660_));
 sky130_fd_sc_hd__nand3_2 _34221_ (.A(_11658_),
    .B(_11659_),
    .C(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__nand3_4 _34222_ (.A(_11654_),
    .B(_11655_),
    .C(_11661_),
    .Y(_11662_));
 sky130_fd_sc_hd__o21ai_2 _34223_ (.A1(_11645_),
    .A2(_11653_),
    .B1(_11660_),
    .Y(_11663_));
 sky130_vsdinv _34224_ (.A(_11263_),
    .Y(_11664_));
 sky130_fd_sc_hd__nand2_1 _34225_ (.A(_11258_),
    .B(_11260_),
    .Y(_11665_));
 sky130_fd_sc_hd__o2bb2ai_4 _34226_ (.A1_N(_11268_),
    .A2_N(_11287_),
    .B1(_11664_),
    .B2(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__nor2_2 _34227_ (.A(_11314_),
    .B(_11312_),
    .Y(_11667_));
 sky130_fd_sc_hd__nor2_8 _34228_ (.A(_11311_),
    .B(_11315_),
    .Y(_11668_));
 sky130_fd_sc_hd__nor2_4 _34229_ (.A(_11667_),
    .B(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__nand3_4 _34230_ (.A(_11658_),
    .B(_11659_),
    .C(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__nand3_4 _34231_ (.A(_11663_),
    .B(_11666_),
    .C(_11670_),
    .Y(_11671_));
 sky130_vsdinv _34232_ (.A(_11271_),
    .Y(_11672_));
 sky130_fd_sc_hd__and2_2 _34233_ (.A(_11272_),
    .B(_11276_),
    .X(_11673_));
 sky130_fd_sc_hd__o2bb2ai_2 _34234_ (.A1_N(_11662_),
    .A2_N(_11671_),
    .B1(_11672_),
    .B2(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__nor2_4 _34235_ (.A(_11673_),
    .B(_11672_),
    .Y(_11675_));
 sky130_fd_sc_hd__nand3_4 _34236_ (.A(_11671_),
    .B(_11662_),
    .C(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__nand2_1 _34237_ (.A(_11674_),
    .B(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand2_1 _34238_ (.A(_11285_),
    .B(_10895_),
    .Y(_11678_));
 sky130_fd_sc_hd__and2_1 _34239_ (.A(_11678_),
    .B(_11292_),
    .X(_11679_));
 sky130_fd_sc_hd__nand2_4 _34240_ (.A(_11677_),
    .B(_11679_),
    .Y(_11680_));
 sky130_fd_sc_hd__nand2_1 _34241_ (.A(_11678_),
    .B(_11292_),
    .Y(_11681_));
 sky130_fd_sc_hd__nand3_4 _34242_ (.A(_11674_),
    .B(_11681_),
    .C(_11676_),
    .Y(_11682_));
 sky130_fd_sc_hd__nand2_4 _34243_ (.A(_11680_),
    .B(_11682_),
    .Y(_11683_));
 sky130_vsdinv _34244_ (.A(_11298_),
    .Y(_11684_));
 sky130_fd_sc_hd__a21oi_4 _34245_ (.A1(_11309_),
    .A2(_11297_),
    .B1(_11684_),
    .Y(_11685_));
 sky130_fd_sc_hd__xor2_4 _34246_ (.A(_11683_),
    .B(_11685_),
    .X(_02652_));
 sky130_fd_sc_hd__a21oi_4 _34247_ (.A1(_11658_),
    .A2(_11669_),
    .B1(_11653_),
    .Y(_11686_));
 sky130_vsdinv _34248_ (.A(_11616_),
    .Y(_11687_));
 sky130_fd_sc_hd__nor2_8 _34249_ (.A(_11687_),
    .B(_11621_),
    .Y(_11688_));
 sky130_vsdinv _34250_ (.A(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__and2_2 _34251_ (.A(_11637_),
    .B(_11636_),
    .X(_11690_));
 sky130_fd_sc_hd__nor2_4 _34252_ (.A(_11689_),
    .B(_11690_),
    .Y(_11691_));
 sky130_fd_sc_hd__and3_2 _34253_ (.A(_11637_),
    .B(_11636_),
    .C(_11689_),
    .X(_11692_));
 sky130_fd_sc_hd__nor2_2 _34254_ (.A(_11514_),
    .B(_11478_),
    .Y(_11693_));
 sky130_fd_sc_hd__nor2_4 _34255_ (.A(_11482_),
    .B(_11693_),
    .Y(_11694_));
 sky130_fd_sc_hd__nand2_2 _34256_ (.A(_19881_),
    .B(_06976_),
    .Y(_11695_));
 sky130_fd_sc_hd__a21o_1 _34257_ (.A1(_06638_),
    .A2(_11061_),
    .B1(_11695_),
    .X(_11696_));
 sky130_fd_sc_hd__nand2_2 _34258_ (.A(_07449_),
    .B(_20118_),
    .Y(_11697_));
 sky130_fd_sc_hd__a21o_1 _34259_ (.A1(_11103_),
    .A2(_10694_),
    .B1(_11697_),
    .X(_11698_));
 sky130_fd_sc_hd__nand2_2 _34260_ (.A(net456),
    .B(_09921_),
    .Y(_11699_));
 sky130_fd_sc_hd__nand3_4 _34261_ (.A(_11696_),
    .B(_11698_),
    .C(_11699_),
    .Y(_11700_));
 sky130_fd_sc_hd__nand3_2 _34262_ (.A(_11463_),
    .B(_06638_),
    .C(_07568_),
    .Y(_11701_));
 sky130_fd_sc_hd__nand2_2 _34263_ (.A(_11695_),
    .B(_11697_),
    .Y(_11702_));
 sky130_fd_sc_hd__o2111ai_4 _34264_ (.A1(_10691_),
    .A2(_11701_),
    .B1(net456),
    .C1(_20115_),
    .D1(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__o21ai_1 _34265_ (.A1(_11411_),
    .A2(_11412_),
    .B1(_11414_),
    .Y(_11704_));
 sky130_fd_sc_hd__nand2_2 _34266_ (.A(_11704_),
    .B(_11415_),
    .Y(_11705_));
 sky130_fd_sc_hd__a21boi_4 _34267_ (.A1(_11700_),
    .A2(_11703_),
    .B1_N(_11705_),
    .Y(_11706_));
 sky130_fd_sc_hd__nor2_1 _34268_ (.A(_11414_),
    .B(_11417_),
    .Y(_11707_));
 sky130_fd_sc_hd__o211a_2 _34269_ (.A1(_11418_),
    .A2(_11707_),
    .B1(_11703_),
    .C1(_11700_),
    .X(_11708_));
 sky130_fd_sc_hd__a21oi_4 _34270_ (.A1(_11464_),
    .A2(_11462_),
    .B1(_11459_),
    .Y(_11709_));
 sky130_fd_sc_hd__o21ai_2 _34271_ (.A1(_11706_),
    .A2(_11708_),
    .B1(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__nand2_2 _34272_ (.A(_11700_),
    .B(_11703_),
    .Y(_11711_));
 sky130_fd_sc_hd__a21oi_4 _34273_ (.A1(_11711_),
    .A2(_11705_),
    .B1(_11709_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand3b_4 _34274_ (.A_N(_11705_),
    .B(_11700_),
    .C(_11703_),
    .Y(_11713_));
 sky130_fd_sc_hd__nand2_1 _34275_ (.A(_11712_),
    .B(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__nand2_1 _34276_ (.A(_11472_),
    .B(_11475_),
    .Y(_11715_));
 sky130_fd_sc_hd__nand2_4 _34277_ (.A(_11715_),
    .B(_11467_),
    .Y(_11716_));
 sky130_fd_sc_hd__nand3_4 _34278_ (.A(_11710_),
    .B(_11714_),
    .C(_11716_),
    .Y(_11717_));
 sky130_fd_sc_hd__o21bai_2 _34279_ (.A1(_11706_),
    .A2(_11708_),
    .B1_N(_11709_),
    .Y(_11718_));
 sky130_fd_sc_hd__nand3b_4 _34280_ (.A_N(_11706_),
    .B(_11713_),
    .C(_11709_),
    .Y(_11719_));
 sky130_fd_sc_hd__nand3b_4 _34281_ (.A_N(_11716_),
    .B(_11718_),
    .C(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__nand3_4 _34282_ (.A(_06357_),
    .B(_06895_),
    .C(_08053_),
    .Y(_11721_));
 sky130_fd_sc_hd__nor2_8 _34283_ (.A(_09732_),
    .B(_11721_),
    .Y(_11722_));
 sky130_fd_sc_hd__clkbuf_4 _34284_ (.A(_08196_),
    .X(_11723_));
 sky130_fd_sc_hd__a22o_1 _34285_ (.A1(_11486_),
    .A2(_11487_),
    .B1(_06208_),
    .B2(_11723_),
    .X(_11724_));
 sky130_fd_sc_hd__nand2_4 _34286_ (.A(_10700_),
    .B(_08450_),
    .Y(_11725_));
 sky130_vsdinv _34287_ (.A(_11725_),
    .Y(_11726_));
 sky130_fd_sc_hd__nand2_1 _34288_ (.A(_11724_),
    .B(_11726_),
    .Y(_11727_));
 sky130_fd_sc_hd__a22oi_4 _34289_ (.A1(_11486_),
    .A2(_11487_),
    .B1(_06208_),
    .B2(_11723_),
    .Y(_11728_));
 sky130_fd_sc_hd__o21ai_2 _34290_ (.A1(_11728_),
    .A2(_11722_),
    .B1(_11725_),
    .Y(_11729_));
 sky130_fd_sc_hd__a21o_1 _34291_ (.A1(_11488_),
    .A2(_11490_),
    .B1(_11485_),
    .X(_11730_));
 sky130_fd_sc_hd__o211ai_4 _34292_ (.A1(_11722_),
    .A2(_11727_),
    .B1(_11729_),
    .C1(_11730_),
    .Y(_11731_));
 sky130_fd_sc_hd__o21ai_4 _34293_ (.A1(_11728_),
    .A2(_11722_),
    .B1(_11726_),
    .Y(_11732_));
 sky130_fd_sc_hd__a21oi_4 _34294_ (.A1(_11488_),
    .A2(_11490_),
    .B1(_11485_),
    .Y(_11733_));
 sky130_fd_sc_hd__buf_6 _34295_ (.A(_09732_),
    .X(_11734_));
 sky130_fd_sc_hd__o211ai_4 _34296_ (.A1(_11734_),
    .A2(_11721_),
    .B1(_11725_),
    .C1(_11724_),
    .Y(_11735_));
 sky130_fd_sc_hd__nand3_4 _34297_ (.A(_11732_),
    .B(_11733_),
    .C(_11735_),
    .Y(_11736_));
 sky130_fd_sc_hd__nand2_8 _34298_ (.A(_11503_),
    .B(_10222_),
    .Y(_11737_));
 sky130_fd_sc_hd__a22o_2 _34299_ (.A1(_06119_),
    .A2(_09044_),
    .B1(_10347_),
    .B2(_09493_),
    .X(_11738_));
 sky130_fd_sc_hd__o21ai_1 _34300_ (.A1(_06623_),
    .A2(_11737_),
    .B1(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__nand2_4 _34301_ (.A(_06052_),
    .B(_09490_),
    .Y(_11740_));
 sky130_vsdinv _34302_ (.A(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__nand2_2 _34303_ (.A(_11739_),
    .B(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__nor2_2 _34304_ (.A(_06623_),
    .B(_11737_),
    .Y(_11743_));
 sky130_fd_sc_hd__nand3b_4 _34305_ (.A_N(_11743_),
    .B(_11740_),
    .C(_11738_),
    .Y(_11744_));
 sky130_fd_sc_hd__nand2_2 _34306_ (.A(_11742_),
    .B(_11744_),
    .Y(_11745_));
 sky130_fd_sc_hd__nand3_2 _34307_ (.A(_11731_),
    .B(_11736_),
    .C(_11745_),
    .Y(_11746_));
 sky130_vsdinv _34308_ (.A(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__nand2_1 _34309_ (.A(_11731_),
    .B(_11736_),
    .Y(_11748_));
 sky130_fd_sc_hd__nand2_1 _34310_ (.A(_11739_),
    .B(_11740_),
    .Y(_11749_));
 sky130_fd_sc_hd__nand3b_2 _34311_ (.A_N(_11743_),
    .B(_11741_),
    .C(_11738_),
    .Y(_11750_));
 sky130_fd_sc_hd__nand2_4 _34312_ (.A(_11749_),
    .B(_11750_),
    .Y(_11751_));
 sky130_fd_sc_hd__nand2_1 _34313_ (.A(_11748_),
    .B(_11751_),
    .Y(_11752_));
 sky130_vsdinv _34314_ (.A(_11752_),
    .Y(_11753_));
 sky130_fd_sc_hd__o2bb2ai_2 _34315_ (.A1_N(_11717_),
    .A2_N(_11720_),
    .B1(_11747_),
    .B2(_11753_),
    .Y(_11754_));
 sky130_fd_sc_hd__and2_1 _34316_ (.A(_11752_),
    .B(_11746_),
    .X(_11755_));
 sky130_fd_sc_hd__nand3_2 _34317_ (.A(_11755_),
    .B(_11717_),
    .C(_11720_),
    .Y(_11756_));
 sky130_fd_sc_hd__o21ai_4 _34318_ (.A1(_11439_),
    .A2(_11440_),
    .B1(_11432_),
    .Y(_11757_));
 sky130_fd_sc_hd__nand3_4 _34319_ (.A(_11754_),
    .B(_11756_),
    .C(_11757_),
    .Y(_11758_));
 sky130_fd_sc_hd__nor2_2 _34320_ (.A(_11745_),
    .B(_11748_),
    .Y(_11759_));
 sky130_vsdinv _34321_ (.A(_11748_),
    .Y(_11760_));
 sky130_fd_sc_hd__nor2_2 _34322_ (.A(_11751_),
    .B(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__o2bb2ai_4 _34323_ (.A1_N(_11717_),
    .A2_N(_11720_),
    .B1(_11759_),
    .B2(_11761_),
    .Y(_11762_));
 sky130_fd_sc_hd__a21oi_4 _34324_ (.A1(_11427_),
    .A2(_11434_),
    .B1(_11450_),
    .Y(_11763_));
 sky130_fd_sc_hd__nand2_1 _34325_ (.A(_11752_),
    .B(_11746_),
    .Y(_11764_));
 sky130_fd_sc_hd__nand3_4 _34326_ (.A(_11720_),
    .B(_11717_),
    .C(_11764_),
    .Y(_11765_));
 sky130_fd_sc_hd__nand3_4 _34327_ (.A(_11762_),
    .B(_11763_),
    .C(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__nand2_1 _34328_ (.A(_11758_),
    .B(_11766_),
    .Y(_11767_));
 sky130_fd_sc_hd__nor2_2 _34329_ (.A(_11694_),
    .B(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__or2_2 _34330_ (.A(_11482_),
    .B(_11693_),
    .X(_11769_));
 sky130_fd_sc_hd__a21oi_4 _34331_ (.A1(_11758_),
    .A2(_11766_),
    .B1(_11769_),
    .Y(_11770_));
 sky130_fd_sc_hd__a21o_1 _34332_ (.A1(_11377_),
    .A2(_11379_),
    .B1(_11381_),
    .X(_11771_));
 sky130_fd_sc_hd__nand2_1 _34333_ (.A(_11387_),
    .B(_11379_),
    .Y(_11772_));
 sky130_fd_sc_hd__nand3_1 _34334_ (.A(_11354_),
    .B(_11771_),
    .C(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand2_2 _34335_ (.A(_11773_),
    .B(_11362_),
    .Y(_11774_));
 sky130_fd_sc_hd__nand3_4 _34336_ (.A(_10961_),
    .B(_10962_),
    .C(_05176_),
    .Y(_11775_));
 sky130_fd_sc_hd__nor2_2 _34337_ (.A(_06197_),
    .B(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__buf_6 _34338_ (.A(\pcpi_mul.rs2[31] ),
    .X(_11777_));
 sky130_fd_sc_hd__buf_4 _34339_ (.A(\pcpi_mul.rs2[32] ),
    .X(_11778_));
 sky130_fd_sc_hd__a22oi_4 _34340_ (.A1(_11777_),
    .A2(_20168_),
    .B1(_05126_),
    .B2(_11778_),
    .Y(_11779_));
 sky130_fd_sc_hd__nand2_4 _34341_ (.A(_19832_),
    .B(_05460_),
    .Y(_11780_));
 sky130_vsdinv _34342_ (.A(_11780_),
    .Y(_11781_));
 sky130_fd_sc_hd__o21ai_2 _34343_ (.A1(_11776_),
    .A2(_11779_),
    .B1(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__buf_6 _34344_ (.A(_10962_),
    .X(_11783_));
 sky130_fd_sc_hd__o2bb2ai_4 _34345_ (.A1_N(_11783_),
    .A2_N(_06614_),
    .B1(_20171_),
    .B2(_10967_),
    .Y(_11784_));
 sky130_fd_sc_hd__o211ai_2 _34346_ (.A1(_05144_),
    .A2(_11775_),
    .B1(_11780_),
    .C1(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__o21ai_1 _34347_ (.A1(_05418_),
    .A2(_11321_),
    .B1(_11324_),
    .Y(_11786_));
 sky130_fd_sc_hd__nand2_1 _34348_ (.A(_11786_),
    .B(_11327_),
    .Y(_11787_));
 sky130_fd_sc_hd__nand3_4 _34349_ (.A(_11782_),
    .B(_11785_),
    .C(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__o21ai_1 _34350_ (.A1(_11776_),
    .A2(_11779_),
    .B1(_11780_),
    .Y(_11789_));
 sky130_fd_sc_hd__o211ai_2 _34351_ (.A1(_20172_),
    .A2(_11775_),
    .B1(_11781_),
    .C1(_11784_),
    .Y(_11790_));
 sky130_fd_sc_hd__o22ai_2 _34352_ (.A1(_05147_),
    .A2(_11321_),
    .B1(_11324_),
    .B2(_11323_),
    .Y(_11791_));
 sky130_fd_sc_hd__nand3_2 _34353_ (.A(_11789_),
    .B(_11790_),
    .C(_11791_),
    .Y(_11792_));
 sky130_fd_sc_hd__buf_2 _34354_ (.A(_11792_),
    .X(_11793_));
 sky130_fd_sc_hd__buf_6 _34355_ (.A(\pcpi_mul.rs2[29] ),
    .X(_11794_));
 sky130_fd_sc_hd__a22oi_4 _34356_ (.A1(_11794_),
    .A2(_05867_),
    .B1(_19840_),
    .B2(_05577_),
    .Y(_11795_));
 sky130_fd_sc_hd__nor2_4 _34357_ (.A(_06624_),
    .B(_10987_),
    .Y(_11796_));
 sky130_fd_sc_hd__nand2_4 _34358_ (.A(_09696_),
    .B(_05696_),
    .Y(_11797_));
 sky130_vsdinv _34359_ (.A(_11797_),
    .Y(_11798_));
 sky130_fd_sc_hd__o21ai_1 _34360_ (.A1(_11795_),
    .A2(_11796_),
    .B1(_11798_),
    .Y(_11799_));
 sky130_vsdinv _34361_ (.A(_11799_),
    .Y(_11800_));
 sky130_fd_sc_hd__or2_1 _34362_ (.A(_06624_),
    .B(_10983_),
    .X(_11801_));
 sky130_fd_sc_hd__a22o_2 _34363_ (.A1(_11794_),
    .A2(_05867_),
    .B1(_19840_),
    .B2(_05577_),
    .X(_11802_));
 sky130_fd_sc_hd__nand3_2 _34364_ (.A(_11801_),
    .B(_11797_),
    .C(_11802_),
    .Y(_11803_));
 sky130_vsdinv _34365_ (.A(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__o2bb2ai_2 _34366_ (.A1_N(_11788_),
    .A2_N(_11793_),
    .B1(_11800_),
    .B2(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__o21ai_1 _34367_ (.A1(_20175_),
    .A2(_11321_),
    .B1(_11327_),
    .Y(_11806_));
 sky130_fd_sc_hd__a21oi_2 _34368_ (.A1(_11806_),
    .A2(_11324_),
    .B1(_11334_),
    .Y(_11807_));
 sky130_fd_sc_hd__a22oi_4 _34369_ (.A1(_11807_),
    .A2(_11328_),
    .B1(_11335_),
    .B2(_11352_),
    .Y(_11808_));
 sky130_fd_sc_hd__o211a_1 _34370_ (.A1(_06624_),
    .A2(_10988_),
    .B1(_11798_),
    .C1(_11802_),
    .X(_11809_));
 sky130_fd_sc_hd__nor2_1 _34371_ (.A(_11795_),
    .B(_11796_),
    .Y(_11810_));
 sky130_fd_sc_hd__nor2_2 _34372_ (.A(_11798_),
    .B(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__o211ai_2 _34373_ (.A1(_11809_),
    .A2(_11811_),
    .B1(_11788_),
    .C1(_11793_),
    .Y(_11812_));
 sky130_fd_sc_hd__nand3_4 _34374_ (.A(_11805_),
    .B(_11808_),
    .C(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__nand2_1 _34375_ (.A(_11335_),
    .B(_11352_),
    .Y(_11814_));
 sky130_fd_sc_hd__nand2_1 _34376_ (.A(_11814_),
    .B(_11330_),
    .Y(_11815_));
 sky130_fd_sc_hd__o2bb2ai_1 _34377_ (.A1_N(_11788_),
    .A2_N(_11793_),
    .B1(_11811_),
    .B2(_11809_),
    .Y(_11816_));
 sky130_fd_sc_hd__nand2_2 _34378_ (.A(_11803_),
    .B(_11799_),
    .Y(_11817_));
 sky130_fd_sc_hd__nand3_1 _34379_ (.A(_11788_),
    .B(_11793_),
    .C(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__nand3_2 _34380_ (.A(_11815_),
    .B(_11816_),
    .C(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__clkbuf_4 _34381_ (.A(_11819_),
    .X(_11820_));
 sky130_fd_sc_hd__nand2_4 _34382_ (.A(_19850_),
    .B(_05827_),
    .Y(_11821_));
 sky130_fd_sc_hd__nand3_2 _34383_ (.A(_11821_),
    .B(_19848_),
    .C(_05979_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand2_4 _34384_ (.A(_19847_),
    .B(_05454_),
    .Y(_11823_));
 sky130_fd_sc_hd__nand3_2 _34385_ (.A(_11823_),
    .B(_11010_),
    .C(_06148_),
    .Y(_11824_));
 sky130_fd_sc_hd__o211ai_4 _34386_ (.A1(_08614_),
    .A2(_06288_),
    .B1(_11822_),
    .C1(_11824_),
    .Y(_11825_));
 sky130_fd_sc_hd__buf_6 _34387_ (.A(_09980_),
    .X(_11826_));
 sky130_fd_sc_hd__nand3_2 _34388_ (.A(_11826_),
    .B(_10384_),
    .C(_06476_),
    .Y(_11827_));
 sky130_fd_sc_hd__and2_1 _34389_ (.A(_19853_),
    .B(_05826_),
    .X(_11828_));
 sky130_fd_sc_hd__nand2_1 _34390_ (.A(_11823_),
    .B(_11821_),
    .Y(_11829_));
 sky130_fd_sc_hd__o211ai_4 _34391_ (.A1(_06672_),
    .A2(_11827_),
    .B1(_11828_),
    .C1(_11829_),
    .Y(_11830_));
 sky130_fd_sc_hd__nand2_1 _34392_ (.A(_11825_),
    .B(_11830_),
    .Y(_11831_));
 sky130_fd_sc_hd__nor2_1 _34393_ (.A(_11345_),
    .B(_11356_),
    .Y(_11832_));
 sky130_fd_sc_hd__nand2_2 _34394_ (.A(_11831_),
    .B(_11832_),
    .Y(_11833_));
 sky130_fd_sc_hd__o2bb2ai_4 _34395_ (.A1_N(_11339_),
    .A2_N(_11342_),
    .B1(_07752_),
    .B2(_11336_),
    .Y(_11834_));
 sky130_fd_sc_hd__nand3_4 _34396_ (.A(_11834_),
    .B(_11825_),
    .C(_11830_),
    .Y(_11835_));
 sky130_fd_sc_hd__nand2_2 _34397_ (.A(_11375_),
    .B(_11372_),
    .Y(_11836_));
 sky130_fd_sc_hd__a21oi_4 _34398_ (.A1(_11833_),
    .A2(_11835_),
    .B1(_11836_),
    .Y(_11837_));
 sky130_fd_sc_hd__a21boi_4 _34399_ (.A1(_11373_),
    .A2(_11374_),
    .B1_N(_11372_),
    .Y(_11838_));
 sky130_fd_sc_hd__a21oi_4 _34400_ (.A1(_11825_),
    .A2(_11830_),
    .B1(_11834_),
    .Y(_11839_));
 sky130_fd_sc_hd__nor2_4 _34401_ (.A(_11838_),
    .B(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__nand2_1 _34402_ (.A(_11840_),
    .B(_11835_),
    .Y(_11841_));
 sky130_vsdinv _34403_ (.A(_11841_),
    .Y(_11842_));
 sky130_fd_sc_hd__o2bb2ai_2 _34404_ (.A1_N(_11813_),
    .A2_N(_11820_),
    .B1(_11837_),
    .B2(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__a21oi_4 _34405_ (.A1(_11835_),
    .A2(_11840_),
    .B1(_11837_),
    .Y(_11844_));
 sky130_fd_sc_hd__nand3_4 _34406_ (.A(_11820_),
    .B(_11813_),
    .C(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__nand3_4 _34407_ (.A(_11774_),
    .B(_11843_),
    .C(_11845_),
    .Y(_11846_));
 sky130_fd_sc_hd__a21o_1 _34408_ (.A1(_11835_),
    .A2(_11840_),
    .B1(_11837_),
    .X(_11847_));
 sky130_fd_sc_hd__a21o_1 _34409_ (.A1(_11820_),
    .A2(_11813_),
    .B1(_11847_),
    .X(_11848_));
 sky130_fd_sc_hd__a21boi_4 _34410_ (.A1(_11388_),
    .A2(_11354_),
    .B1_N(_11362_),
    .Y(_11849_));
 sky130_fd_sc_hd__nand3_2 _34411_ (.A(_11847_),
    .B(_11820_),
    .C(_11813_),
    .Y(_11850_));
 sky130_fd_sc_hd__nand3_4 _34412_ (.A(_11848_),
    .B(_11849_),
    .C(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__nand3_4 _34413_ (.A(_19858_),
    .B(_08575_),
    .C(_07024_),
    .Y(_11852_));
 sky130_fd_sc_hd__nor2_8 _34414_ (.A(net465),
    .B(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__a22o_2 _34415_ (.A1(_10433_),
    .A2(_06154_),
    .B1(_10620_),
    .B2(_06151_),
    .X(_11854_));
 sky130_fd_sc_hd__nand2_4 _34416_ (.A(_10435_),
    .B(_07661_),
    .Y(_11855_));
 sky130_vsdinv _34417_ (.A(_11855_),
    .Y(_11856_));
 sky130_fd_sc_hd__nand2_1 _34418_ (.A(_11854_),
    .B(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__o22ai_4 _34419_ (.A1(_06308_),
    .A2(_11398_),
    .B1(_11400_),
    .B2(_11397_),
    .Y(_11858_));
 sky130_fd_sc_hd__a22oi_4 _34420_ (.A1(_10433_),
    .A2(_06154_),
    .B1(_10620_),
    .B2(_06151_),
    .Y(_11859_));
 sky130_fd_sc_hd__o21ai_2 _34421_ (.A1(_11859_),
    .A2(_11853_),
    .B1(_11855_),
    .Y(_11860_));
 sky130_fd_sc_hd__o211ai_4 _34422_ (.A1(_11853_),
    .A2(_11857_),
    .B1(_11858_),
    .C1(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__o21ai_2 _34423_ (.A1(_11859_),
    .A2(_11853_),
    .B1(_11856_),
    .Y(_11862_));
 sky130_fd_sc_hd__a21oi_2 _34424_ (.A1(_11404_),
    .A2(_11401_),
    .B1(_11399_),
    .Y(_11863_));
 sky130_fd_sc_hd__o211ai_4 _34425_ (.A1(_07191_),
    .A2(_11852_),
    .B1(_11855_),
    .C1(_11854_),
    .Y(_11864_));
 sky130_fd_sc_hd__nand3_4 _34426_ (.A(_11862_),
    .B(_11863_),
    .C(_11864_),
    .Y(_11865_));
 sky130_fd_sc_hd__nand2_1 _34427_ (.A(_11861_),
    .B(_11865_),
    .Y(_11866_));
 sky130_fd_sc_hd__nand2_1 _34428_ (.A(_19870_),
    .B(_08546_),
    .Y(_11867_));
 sky130_fd_sc_hd__nand3b_2 _34429_ (.A_N(_11867_),
    .B(_10945_),
    .C(_20131_),
    .Y(_11868_));
 sky130_fd_sc_hd__buf_4 _34430_ (.A(_19876_),
    .X(_11869_));
 sky130_fd_sc_hd__nand2_4 _34431_ (.A(_11869_),
    .B(_07258_),
    .Y(_11870_));
 sky130_fd_sc_hd__buf_4 _34432_ (.A(_19873_),
    .X(_11871_));
 sky130_fd_sc_hd__nand2_1 _34433_ (.A(_11871_),
    .B(_11093_),
    .Y(_11872_));
 sky130_fd_sc_hd__nand2_1 _34434_ (.A(_11867_),
    .B(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__and3_2 _34435_ (.A(_11868_),
    .B(_11870_),
    .C(_11873_),
    .X(_11874_));
 sky130_fd_sc_hd__a22oi_4 _34436_ (.A1(_10935_),
    .A2(_20134_),
    .B1(_10945_),
    .B2(_20131_),
    .Y(_11875_));
 sky130_fd_sc_hd__nor2_1 _34437_ (.A(_11867_),
    .B(_11872_),
    .Y(_11876_));
 sky130_fd_sc_hd__nor2_2 _34438_ (.A(_11875_),
    .B(_11876_),
    .Y(_11877_));
 sky130_fd_sc_hd__nor2_4 _34439_ (.A(_11870_),
    .B(_11877_),
    .Y(_11878_));
 sky130_fd_sc_hd__nor2_8 _34440_ (.A(_11874_),
    .B(_11878_),
    .Y(_11879_));
 sky130_fd_sc_hd__nand2_4 _34441_ (.A(_11866_),
    .B(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__a21o_1 _34442_ (.A1(_11868_),
    .A2(_11873_),
    .B1(_11870_),
    .X(_11881_));
 sky130_fd_sc_hd__nand2_1 _34443_ (.A(_11877_),
    .B(_11870_),
    .Y(_11882_));
 sky130_fd_sc_hd__nand2_4 _34444_ (.A(_11881_),
    .B(_11882_),
    .Y(_11883_));
 sky130_fd_sc_hd__nand3_4 _34445_ (.A(_11883_),
    .B(_11865_),
    .C(_11861_),
    .Y(_11884_));
 sky130_fd_sc_hd__a21oi_4 _34446_ (.A1(_11380_),
    .A2(_11379_),
    .B1(_11386_),
    .Y(_11885_));
 sky130_fd_sc_hd__a21o_2 _34447_ (.A1(_11880_),
    .A2(_11884_),
    .B1(_11885_),
    .X(_11886_));
 sky130_fd_sc_hd__nand3_4 _34448_ (.A(_11880_),
    .B(_11885_),
    .C(_11884_),
    .Y(_11887_));
 sky130_fd_sc_hd__nand2_4 _34449_ (.A(_11431_),
    .B(_11410_),
    .Y(_11888_));
 sky130_fd_sc_hd__a21oi_2 _34450_ (.A1(_11886_),
    .A2(_11887_),
    .B1(_11888_),
    .Y(_11889_));
 sky130_fd_sc_hd__and3_1 _34451_ (.A(_11886_),
    .B(_11888_),
    .C(_11887_),
    .X(_11890_));
 sky130_fd_sc_hd__o2bb2ai_4 _34452_ (.A1_N(_11846_),
    .A2_N(_11851_),
    .B1(_11889_),
    .B2(_11890_),
    .Y(_11891_));
 sky130_fd_sc_hd__a21oi_4 _34453_ (.A1(_11880_),
    .A2(_11884_),
    .B1(_11885_),
    .Y(_11892_));
 sky130_fd_sc_hd__and3_2 _34454_ (.A(_11880_),
    .B(_11885_),
    .C(_11884_),
    .X(_11893_));
 sky130_fd_sc_hd__o21ai_2 _34455_ (.A1(_11892_),
    .A2(_11893_),
    .B1(_11888_),
    .Y(_11894_));
 sky130_fd_sc_hd__and2_2 _34456_ (.A(_11431_),
    .B(_11410_),
    .X(_11895_));
 sky130_fd_sc_hd__nand3_2 _34457_ (.A(_11886_),
    .B(_11895_),
    .C(_11887_),
    .Y(_11896_));
 sky130_fd_sc_hd__nand2_4 _34458_ (.A(_11894_),
    .B(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__nand3_4 _34459_ (.A(_11897_),
    .B(_11851_),
    .C(_11846_),
    .Y(_11898_));
 sky130_fd_sc_hd__nand2_1 _34460_ (.A(_11442_),
    .B(_11395_),
    .Y(_11899_));
 sky130_fd_sc_hd__nand2_2 _34461_ (.A(_11899_),
    .B(_11390_),
    .Y(_11900_));
 sky130_fd_sc_hd__a21oi_4 _34462_ (.A1(_11891_),
    .A2(_11898_),
    .B1(_11900_),
    .Y(_11901_));
 sky130_vsdinv _34463_ (.A(_11390_),
    .Y(_11902_));
 sky130_fd_sc_hd__nand2_1 _34464_ (.A(_11384_),
    .B(_11389_),
    .Y(_11903_));
 sky130_fd_sc_hd__a21oi_4 _34465_ (.A1(_11903_),
    .A2(_11393_),
    .B1(_11452_),
    .Y(_11904_));
 sky130_fd_sc_hd__o211a_2 _34466_ (.A1(_11902_),
    .A2(_11904_),
    .B1(_11898_),
    .C1(_11891_),
    .X(_11905_));
 sky130_fd_sc_hd__o22ai_4 _34467_ (.A1(_11768_),
    .A2(_11770_),
    .B1(_11901_),
    .B2(_11905_),
    .Y(_11906_));
 sky130_fd_sc_hd__a21oi_2 _34468_ (.A1(_11851_),
    .A2(_11846_),
    .B1(_11897_),
    .Y(_11907_));
 sky130_fd_sc_hd__a21oi_1 _34469_ (.A1(_11886_),
    .A2(_11887_),
    .B1(_11895_),
    .Y(_11908_));
 sky130_fd_sc_hd__nor3_2 _34470_ (.A(_11888_),
    .B(_11892_),
    .C(_11893_),
    .Y(_11909_));
 sky130_fd_sc_hd__o211a_1 _34471_ (.A1(_11908_),
    .A2(_11909_),
    .B1(_11846_),
    .C1(_11851_),
    .X(_11910_));
 sky130_fd_sc_hd__nor2_2 _34472_ (.A(_11902_),
    .B(_11904_),
    .Y(_11911_));
 sky130_fd_sc_hd__o21ai_4 _34473_ (.A1(_11907_),
    .A2(_11910_),
    .B1(_11911_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand3_4 _34474_ (.A(_11900_),
    .B(_11898_),
    .C(_11891_),
    .Y(_11913_));
 sky130_fd_sc_hd__a31oi_4 _34475_ (.A1(_11763_),
    .A2(_11762_),
    .A3(_11765_),
    .B1(_11694_),
    .Y(_11914_));
 sky130_fd_sc_hd__a21oi_4 _34476_ (.A1(_11758_),
    .A2(_11914_),
    .B1(_11770_),
    .Y(_11915_));
 sky130_fd_sc_hd__nand3_4 _34477_ (.A(_11912_),
    .B(_11913_),
    .C(_11915_),
    .Y(_11916_));
 sky130_fd_sc_hd__a21oi_2 _34478_ (.A1(_11438_),
    .A2(_11443_),
    .B1(_11320_),
    .Y(_11917_));
 sky130_fd_sc_hd__o21ai_4 _34479_ (.A1(_11541_),
    .A2(_11917_),
    .B1(_11444_),
    .Y(_11918_));
 sky130_fd_sc_hd__nand3_4 _34480_ (.A(_11906_),
    .B(_11916_),
    .C(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__o21ai_2 _34481_ (.A1(_11901_),
    .A2(_11905_),
    .B1(_11915_),
    .Y(_11920_));
 sky130_fd_sc_hd__a21boi_4 _34482_ (.A1(_11533_),
    .A2(_11454_),
    .B1_N(_11444_),
    .Y(_11921_));
 sky130_fd_sc_hd__nand2_1 _34483_ (.A(_11914_),
    .B(_11758_),
    .Y(_11922_));
 sky130_fd_sc_hd__nand2_1 _34484_ (.A(_11767_),
    .B(_11694_),
    .Y(_11923_));
 sky130_fd_sc_hd__nand2_2 _34485_ (.A(_11922_),
    .B(_11923_),
    .Y(_11924_));
 sky130_fd_sc_hd__nand3_4 _34486_ (.A(_11912_),
    .B(_11913_),
    .C(_11924_),
    .Y(_11925_));
 sky130_fd_sc_hd__nand3_4 _34487_ (.A(_11920_),
    .B(_11921_),
    .C(_11925_),
    .Y(_11926_));
 sky130_fd_sc_hd__buf_4 _34488_ (.A(_09025_),
    .X(_11927_));
 sky130_fd_sc_hd__a22oi_4 _34489_ (.A1(_19913_),
    .A2(_11927_),
    .B1(_19916_),
    .B2(_10262_),
    .Y(_11928_));
 sky130_fd_sc_hd__nand3_4 _34490_ (.A(_05858_),
    .B(_05414_),
    .C(_20086_),
    .Y(_11929_));
 sky130_fd_sc_hd__nor2_2 _34491_ (.A(_10781_),
    .B(_11929_),
    .Y(_11930_));
 sky130_fd_sc_hd__nand2_2 _34492_ (.A(_05866_),
    .B(_09896_),
    .Y(_11931_));
 sky130_fd_sc_hd__o21ai_2 _34493_ (.A1(_11928_),
    .A2(_11930_),
    .B1(_11931_),
    .Y(_11932_));
 sky130_vsdinv _34494_ (.A(_11931_),
    .Y(_11933_));
 sky130_fd_sc_hd__buf_4 _34495_ (.A(_20085_),
    .X(_11934_));
 sky130_fd_sc_hd__a22o_1 _34496_ (.A1(_10809_),
    .A2(_20091_),
    .B1(_11206_),
    .B2(_11934_),
    .X(_11935_));
 sky130_fd_sc_hd__o211ai_2 _34497_ (.A1(_10781_),
    .A2(_11929_),
    .B1(_11933_),
    .C1(_11935_),
    .Y(_11936_));
 sky130_fd_sc_hd__o21ai_2 _34498_ (.A1(_11504_),
    .A2(_11501_),
    .B1(_11508_),
    .Y(_11937_));
 sky130_fd_sc_hd__nand3_4 _34499_ (.A(_11932_),
    .B(_11936_),
    .C(_11937_),
    .Y(_11938_));
 sky130_fd_sc_hd__o21ai_2 _34500_ (.A1(_11928_),
    .A2(_11930_),
    .B1(_11933_),
    .Y(_11939_));
 sky130_fd_sc_hd__a21oi_4 _34501_ (.A1(_11509_),
    .A2(_11505_),
    .B1(_11502_),
    .Y(_11940_));
 sky130_fd_sc_hd__buf_6 _34502_ (.A(_10780_),
    .X(_11941_));
 sky130_fd_sc_hd__o211ai_2 _34503_ (.A1(_11941_),
    .A2(_11929_),
    .B1(_11931_),
    .C1(_11935_),
    .Y(_11942_));
 sky130_fd_sc_hd__nand3_4 _34504_ (.A(_11939_),
    .B(_11940_),
    .C(_11942_),
    .Y(_11943_));
 sky130_fd_sc_hd__nor2_8 _34505_ (.A(_11553_),
    .B(_11551_),
    .Y(_11944_));
 sky130_fd_sc_hd__o2bb2ai_4 _34506_ (.A1_N(_11938_),
    .A2_N(_11943_),
    .B1(_11548_),
    .B2(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__nor2_4 _34507_ (.A(_11548_),
    .B(_11944_),
    .Y(_11946_));
 sky130_fd_sc_hd__nand3_4 _34508_ (.A(_11943_),
    .B(_11938_),
    .C(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__nand2_4 _34509_ (.A(_11512_),
    .B(_11495_),
    .Y(_11948_));
 sky130_fd_sc_hd__a21oi_4 _34510_ (.A1(_11945_),
    .A2(_11947_),
    .B1(_11948_),
    .Y(_11949_));
 sky130_fd_sc_hd__and3_1 _34511_ (.A(_11948_),
    .B(_11945_),
    .C(_11947_),
    .X(_11950_));
 sky130_fd_sc_hd__nand2_2 _34512_ (.A(_11573_),
    .B(_11565_),
    .Y(_11951_));
 sky130_fd_sc_hd__o21ai_2 _34513_ (.A1(_11949_),
    .A2(_11950_),
    .B1(_11951_),
    .Y(_11952_));
 sky130_fd_sc_hd__a21oi_4 _34514_ (.A1(_11576_),
    .A2(_11578_),
    .B1(_11574_),
    .Y(_11953_));
 sky130_vsdinv _34515_ (.A(_11951_),
    .Y(_11954_));
 sky130_fd_sc_hd__nand3_4 _34516_ (.A(_11948_),
    .B(_11945_),
    .C(_11947_),
    .Y(_11955_));
 sky130_fd_sc_hd__nand3b_4 _34517_ (.A_N(_11949_),
    .B(_11954_),
    .C(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__nand3_4 _34518_ (.A(_11952_),
    .B(_11953_),
    .C(_11956_),
    .Y(_11957_));
 sky130_fd_sc_hd__o21ai_2 _34519_ (.A1(_11949_),
    .A2(_11950_),
    .B1(_11954_),
    .Y(_11958_));
 sky130_fd_sc_hd__o21ai_2 _34520_ (.A1(_11579_),
    .A2(_11571_),
    .B1(_11577_),
    .Y(_11959_));
 sky130_fd_sc_hd__nand3b_2 _34521_ (.A_N(_11949_),
    .B(_11951_),
    .C(_11955_),
    .Y(_11960_));
 sky130_fd_sc_hd__nand3_4 _34522_ (.A(_11958_),
    .B(_11959_),
    .C(_11960_),
    .Y(_11961_));
 sky130_fd_sc_hd__a22oi_4 _34523_ (.A1(_05229_),
    .A2(_20078_),
    .B1(_05805_),
    .B2(_10760_),
    .Y(_11962_));
 sky130_fd_sc_hd__and4_4 _34524_ (.A(_05228_),
    .B(_06988_),
    .C(\pcpi_mul.rs1[30] ),
    .D(_20077_),
    .X(_11963_));
 sky130_fd_sc_hd__clkbuf_4 _34525_ (.A(_11963_),
    .X(_11964_));
 sky130_fd_sc_hd__a211o_1 _34526_ (.A1(_18687_),
    .A2(_19939_),
    .B1(_11962_),
    .C1(_11964_),
    .X(_11965_));
 sky130_fd_sc_hd__nor2_2 _34527_ (.A(_11595_),
    .B(_11589_),
    .Y(_11966_));
 sky130_fd_sc_hd__o21ai_2 _34528_ (.A1(_11962_),
    .A2(_11964_),
    .B1(_11162_),
    .Y(_11967_));
 sky130_fd_sc_hd__nand3_4 _34529_ (.A(_11965_),
    .B(_11966_),
    .C(_11967_),
    .Y(_11968_));
 sky130_fd_sc_hd__a22o_1 _34530_ (.A1(_19921_),
    .A2(_10761_),
    .B1(_19926_),
    .B2(_11174_),
    .X(_11969_));
 sky130_fd_sc_hd__nand2_1 _34531_ (.A(_11969_),
    .B(_11162_),
    .Y(_11970_));
 sky130_fd_sc_hd__o21ai_2 _34532_ (.A1(_11962_),
    .A2(_11964_),
    .B1(_11168_),
    .Y(_11971_));
 sky130_fd_sc_hd__o221ai_4 _34533_ (.A1(_11595_),
    .A2(_11589_),
    .B1(_11964_),
    .B2(_11970_),
    .C1(_11971_),
    .Y(_11972_));
 sky130_fd_sc_hd__nand2_2 _34534_ (.A(_19928_),
    .B(_20070_),
    .Y(_11973_));
 sky130_fd_sc_hd__o21a_4 _34535_ (.A1(_05387_),
    .A2(_05570_),
    .B1(_18685_),
    .X(_11974_));
 sky130_fd_sc_hd__clkbuf_2 _34536_ (.A(\pcpi_mul.rs1[32] ),
    .X(_11975_));
 sky130_fd_sc_hd__nand3_4 _34537_ (.A(net504),
    .B(_05139_),
    .C(_05477_),
    .Y(_11976_));
 sky130_fd_sc_hd__nand2_2 _34538_ (.A(_11974_),
    .B(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__xor2_4 _34539_ (.A(_11973_),
    .B(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__a21o_1 _34540_ (.A1(_11968_),
    .A2(_11972_),
    .B1(_11978_),
    .X(_11979_));
 sky130_fd_sc_hd__nand3_4 _34541_ (.A(_11978_),
    .B(_11968_),
    .C(_11972_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_1 _34542_ (.A(_11612_),
    .B(_11602_),
    .Y(_11981_));
 sky130_fd_sc_hd__nand2_2 _34543_ (.A(_11981_),
    .B(_11597_),
    .Y(_11982_));
 sky130_fd_sc_hd__a21o_1 _34544_ (.A1(_11979_),
    .A2(_11980_),
    .B1(_11982_),
    .X(_11983_));
 sky130_fd_sc_hd__nand3_2 _34545_ (.A(_11979_),
    .B(_11982_),
    .C(_11980_),
    .Y(_11984_));
 sky130_fd_sc_hd__nor2_4 _34546_ (.A(_11606_),
    .B(_11610_),
    .Y(_11985_));
 sky130_vsdinv _34547_ (.A(_11985_),
    .Y(_11986_));
 sky130_fd_sc_hd__and3_1 _34548_ (.A(_11983_),
    .B(_11984_),
    .C(_11986_),
    .X(_11987_));
 sky130_fd_sc_hd__a21oi_1 _34549_ (.A1(_11983_),
    .A2(_11984_),
    .B1(_11986_),
    .Y(_11988_));
 sky130_fd_sc_hd__o2bb2ai_2 _34550_ (.A1_N(_11957_),
    .A2_N(_11961_),
    .B1(_11987_),
    .B2(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__a21oi_4 _34551_ (.A1(_11979_),
    .A2(_11980_),
    .B1(_11982_),
    .Y(_11990_));
 sky130_fd_sc_hd__and3_1 _34552_ (.A(_11979_),
    .B(_11982_),
    .C(_11980_),
    .X(_11991_));
 sky130_fd_sc_hd__o21ai_1 _34553_ (.A1(_11990_),
    .A2(_11991_),
    .B1(_11986_),
    .Y(_11992_));
 sky130_fd_sc_hd__nand3_1 _34554_ (.A(_11983_),
    .B(_11984_),
    .C(_11985_),
    .Y(_11993_));
 sky130_fd_sc_hd__nand2_2 _34555_ (.A(_11992_),
    .B(_11993_),
    .Y(_11994_));
 sky130_fd_sc_hd__nand3_4 _34556_ (.A(_11994_),
    .B(_11957_),
    .C(_11961_),
    .Y(_11995_));
 sky130_fd_sc_hd__nand2_2 _34557_ (.A(_11529_),
    .B(_11530_),
    .Y(_11996_));
 sky130_fd_sc_hd__nand2_1 _34558_ (.A(_11996_),
    .B(_11526_),
    .Y(_11997_));
 sky130_fd_sc_hd__a21o_1 _34559_ (.A1(_11989_),
    .A2(_11995_),
    .B1(_11997_),
    .X(_11998_));
 sky130_fd_sc_hd__nand2_1 _34560_ (.A(_11961_),
    .B(_11957_),
    .Y(_11999_));
 sky130_fd_sc_hd__nor2_2 _34561_ (.A(_11985_),
    .B(_11990_),
    .Y(_12000_));
 sky130_fd_sc_hd__nand2_1 _34562_ (.A(_12000_),
    .B(_11984_),
    .Y(_12001_));
 sky130_fd_sc_hd__o21ai_1 _34563_ (.A1(_11990_),
    .A2(_11991_),
    .B1(_11985_),
    .Y(_12002_));
 sky130_fd_sc_hd__nand2_2 _34564_ (.A(_12001_),
    .B(_12002_),
    .Y(_12003_));
 sky130_fd_sc_hd__a22oi_4 _34565_ (.A1(_11996_),
    .A2(_11526_),
    .B1(_11999_),
    .B2(_12003_),
    .Y(_12004_));
 sky130_fd_sc_hd__nand2_4 _34566_ (.A(_12004_),
    .B(_11995_),
    .Y(_12005_));
 sky130_vsdinv _34567_ (.A(_11581_),
    .Y(_12006_));
 sky130_fd_sc_hd__o21ai_2 _34568_ (.A1(_11630_),
    .A2(_12006_),
    .B1(_11586_),
    .Y(_12007_));
 sky130_fd_sc_hd__a21oi_2 _34569_ (.A1(_11998_),
    .A2(_12005_),
    .B1(_12007_),
    .Y(_12008_));
 sky130_fd_sc_hd__and3_1 _34570_ (.A(_11989_),
    .B(_11997_),
    .C(_11995_),
    .X(_12009_));
 sky130_fd_sc_hd__nand2_2 _34571_ (.A(_11998_),
    .B(_12007_),
    .Y(_12010_));
 sky130_fd_sc_hd__nor2_2 _34572_ (.A(_12009_),
    .B(_12010_),
    .Y(_12011_));
 sky130_fd_sc_hd__o2bb2ai_4 _34573_ (.A1_N(_11919_),
    .A2_N(_11926_),
    .B1(_12008_),
    .B2(_12011_),
    .Y(_12012_));
 sky130_vsdinv _34574_ (.A(_11586_),
    .Y(_12013_));
 sky130_fd_sc_hd__nor2_2 _34575_ (.A(_11630_),
    .B(_12006_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21oi_2 _34576_ (.A1(_11989_),
    .A2(_11995_),
    .B1(_11997_),
    .Y(_12015_));
 sky130_fd_sc_hd__o22ai_4 _34577_ (.A1(_12013_),
    .A2(_12014_),
    .B1(_12015_),
    .B2(_12009_),
    .Y(_12016_));
 sky130_vsdinv _34578_ (.A(_12007_),
    .Y(_12017_));
 sky130_fd_sc_hd__nand3_4 _34579_ (.A(_11998_),
    .B(_12005_),
    .C(_12017_),
    .Y(_12018_));
 sky130_fd_sc_hd__nand2_4 _34580_ (.A(_12016_),
    .B(_12018_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand3_4 _34581_ (.A(_12019_),
    .B(_11926_),
    .C(_11919_),
    .Y(_12020_));
 sky130_fd_sc_hd__a21oi_2 _34582_ (.A1(_11532_),
    .A2(_11534_),
    .B1(_11317_),
    .Y(_12021_));
 sky130_fd_sc_hd__o21ai_4 _34583_ (.A1(_11649_),
    .A2(_12021_),
    .B1(_11536_),
    .Y(_12022_));
 sky130_fd_sc_hd__a21oi_4 _34584_ (.A1(_12012_),
    .A2(_12020_),
    .B1(_12022_),
    .Y(_12023_));
 sky130_fd_sc_hd__and3_1 _34585_ (.A(_11906_),
    .B(_11918_),
    .C(_11916_),
    .X(_12024_));
 sky130_fd_sc_hd__nand2_2 _34586_ (.A(_12019_),
    .B(_11926_),
    .Y(_12025_));
 sky130_fd_sc_hd__o211a_2 _34587_ (.A1(_12024_),
    .A2(_12025_),
    .B1(_12022_),
    .C1(_12012_),
    .X(_12026_));
 sky130_fd_sc_hd__o22ai_4 _34588_ (.A1(_11691_),
    .A2(_11692_),
    .B1(_12023_),
    .B2(_12026_),
    .Y(_12027_));
 sky130_fd_sc_hd__a21oi_4 _34589_ (.A1(_11926_),
    .A2(_11919_),
    .B1(_12019_),
    .Y(_12028_));
 sky130_fd_sc_hd__a21oi_1 _34590_ (.A1(_11912_),
    .A2(_11913_),
    .B1(_11915_),
    .Y(_12029_));
 sky130_fd_sc_hd__nand2_1 _34591_ (.A(_11918_),
    .B(_11916_),
    .Y(_12030_));
 sky130_fd_sc_hd__o211a_1 _34592_ (.A1(_12029_),
    .A2(_12030_),
    .B1(_11926_),
    .C1(_12019_),
    .X(_12031_));
 sky130_fd_sc_hd__o21bai_4 _34593_ (.A1(_12028_),
    .A2(_12031_),
    .B1_N(_12022_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand3_4 _34594_ (.A(_12012_),
    .B(_12022_),
    .C(_12020_),
    .Y(_12033_));
 sky130_fd_sc_hd__nor2_4 _34595_ (.A(_11692_),
    .B(_11691_),
    .Y(_12034_));
 sky130_fd_sc_hd__nand3_4 _34596_ (.A(_12032_),
    .B(_12033_),
    .C(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__nand3_4 _34597_ (.A(_11686_),
    .B(_12027_),
    .C(_12035_),
    .Y(_12036_));
 sky130_fd_sc_hd__nor2_8 _34598_ (.A(_11688_),
    .B(_11690_),
    .Y(_12037_));
 sky130_fd_sc_hd__and3_2 _34599_ (.A(_11637_),
    .B(_11636_),
    .C(_11688_),
    .X(_12038_));
 sky130_fd_sc_hd__o22ai_4 _34600_ (.A1(_12037_),
    .A2(_12038_),
    .B1(_12023_),
    .B2(_12026_),
    .Y(_12039_));
 sky130_fd_sc_hd__o21ai_2 _34601_ (.A1(_11660_),
    .A2(_11645_),
    .B1(_11659_),
    .Y(_12040_));
 sky130_fd_sc_hd__nor2_4 _34602_ (.A(_12038_),
    .B(_12037_),
    .Y(_12041_));
 sky130_fd_sc_hd__nand3_4 _34603_ (.A(_12032_),
    .B(_12033_),
    .C(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__nand3_4 _34604_ (.A(_12039_),
    .B(_12040_),
    .C(_12042_),
    .Y(_12043_));
 sky130_fd_sc_hd__nand3_4 _34605_ (.A(_12036_),
    .B(_12043_),
    .C(_11668_),
    .Y(_12044_));
 sky130_fd_sc_hd__o2bb2ai_2 _34606_ (.A1_N(_12043_),
    .A2_N(_12036_),
    .B1(_11311_),
    .B2(_11315_),
    .Y(_12045_));
 sky130_vsdinv _34607_ (.A(_11662_),
    .Y(_12046_));
 sky130_fd_sc_hd__o21a_4 _34608_ (.A1(_11672_),
    .A2(_11673_),
    .B1(_11671_),
    .X(_12047_));
 sky130_fd_sc_hd__o2bb2ai_2 _34609_ (.A1_N(_12044_),
    .A2_N(_12045_),
    .B1(_12046_),
    .B2(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__nand2_2 _34610_ (.A(_11662_),
    .B(_11675_),
    .Y(_12049_));
 sky130_fd_sc_hd__nand2_8 _34611_ (.A(_12049_),
    .B(_11671_),
    .Y(_12050_));
 sky130_fd_sc_hd__nand3_4 _34612_ (.A(_12050_),
    .B(_12045_),
    .C(_12044_),
    .Y(_12051_));
 sky130_fd_sc_hd__and2_2 _34613_ (.A(_12048_),
    .B(_12051_),
    .X(_12052_));
 sky130_fd_sc_hd__nor2_8 _34614_ (.A(_11299_),
    .B(_11683_),
    .Y(_12053_));
 sky130_fd_sc_hd__nand2_2 _34615_ (.A(_11682_),
    .B(_11298_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand2_8 _34616_ (.A(_12054_),
    .B(_11680_),
    .Y(_12055_));
 sky130_fd_sc_hd__a21boi_4 _34617_ (.A1(net409),
    .A2(_12053_),
    .B1_N(_12055_),
    .Y(_12056_));
 sky130_fd_sc_hd__xnor2_4 _34618_ (.A(_12052_),
    .B(_12056_),
    .Y(_02653_));
 sky130_fd_sc_hd__and2_1 _34619_ (.A(_11887_),
    .B(_11895_),
    .X(_12057_));
 sky130_fd_sc_hd__o21a_1 _34620_ (.A1(_11705_),
    .A2(_11711_),
    .B1(_11709_),
    .X(_12058_));
 sky130_fd_sc_hd__buf_4 _34621_ (.A(_06993_),
    .X(_12059_));
 sky130_fd_sc_hd__a22oi_4 _34622_ (.A1(_11103_),
    .A2(_12059_),
    .B1(_11094_),
    .B2(_10113_),
    .Y(_12060_));
 sky130_fd_sc_hd__nand3_4 _34623_ (.A(_07446_),
    .B(_19886_),
    .C(_08042_),
    .Y(_12061_));
 sky130_fd_sc_hd__nor2_8 _34624_ (.A(_11057_),
    .B(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_2 _34625_ (.A(_06640_),
    .B(_07548_),
    .Y(_12063_));
 sky130_fd_sc_hd__o21ai_2 _34626_ (.A1(_12060_),
    .A2(_12062_),
    .B1(_12063_),
    .Y(_12064_));
 sky130_vsdinv _34627_ (.A(_12063_),
    .Y(_12065_));
 sky130_fd_sc_hd__a22o_2 _34628_ (.A1(_11463_),
    .A2(_11061_),
    .B1(_06638_),
    .B2(_11062_),
    .X(_12066_));
 sky130_fd_sc_hd__o211ai_4 _34629_ (.A1(_11074_),
    .A2(_12061_),
    .B1(_12065_),
    .C1(_12066_),
    .Y(_12067_));
 sky130_fd_sc_hd__o21ai_2 _34630_ (.A1(_11870_),
    .A2(_11875_),
    .B1(_11868_),
    .Y(_12068_));
 sky130_fd_sc_hd__nand3_4 _34631_ (.A(_12064_),
    .B(_12067_),
    .C(_12068_),
    .Y(_12069_));
 sky130_fd_sc_hd__o21ai_2 _34632_ (.A1(_12060_),
    .A2(_12062_),
    .B1(_12065_),
    .Y(_12070_));
 sky130_fd_sc_hd__o21ai_1 _34633_ (.A1(_11867_),
    .A2(_11872_),
    .B1(_11870_),
    .Y(_12071_));
 sky130_fd_sc_hd__nand2_1 _34634_ (.A(_12071_),
    .B(_11873_),
    .Y(_12072_));
 sky130_fd_sc_hd__buf_6 _34635_ (.A(_09602_),
    .X(_12073_));
 sky130_fd_sc_hd__o211ai_4 _34636_ (.A1(_12073_),
    .A2(_12061_),
    .B1(_12063_),
    .C1(_12066_),
    .Y(_12074_));
 sky130_fd_sc_hd__nand3_4 _34637_ (.A(_12070_),
    .B(_12072_),
    .C(_12074_),
    .Y(_12075_));
 sky130_fd_sc_hd__nor2_2 _34638_ (.A(_11695_),
    .B(_11697_),
    .Y(_12076_));
 sky130_fd_sc_hd__a31o_4 _34639_ (.A1(_11702_),
    .A2(net456),
    .A3(_20116_),
    .B1(_12076_),
    .X(_12077_));
 sky130_fd_sc_hd__a21oi_2 _34640_ (.A1(_12069_),
    .A2(_12075_),
    .B1(_12077_),
    .Y(_12078_));
 sky130_fd_sc_hd__a21oi_2 _34641_ (.A1(_11696_),
    .A2(_11698_),
    .B1(_11699_),
    .Y(_12079_));
 sky130_fd_sc_hd__o211a_4 _34642_ (.A1(_12076_),
    .A2(_12079_),
    .B1(_12069_),
    .C1(_12075_),
    .X(_12080_));
 sky130_fd_sc_hd__o22ai_4 _34643_ (.A1(_11706_),
    .A2(_12058_),
    .B1(_12078_),
    .B2(_12080_),
    .Y(_12081_));
 sky130_fd_sc_hd__nand3_2 _34644_ (.A(_12069_),
    .B(_12075_),
    .C(_12077_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_1 _34645_ (.A(_12069_),
    .B(_12075_),
    .Y(_12083_));
 sky130_vsdinv _34646_ (.A(_12077_),
    .Y(_12084_));
 sky130_fd_sc_hd__nand2_1 _34647_ (.A(_12083_),
    .B(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__o211ai_4 _34648_ (.A1(_11708_),
    .A2(_11712_),
    .B1(_12082_),
    .C1(_12085_),
    .Y(_12086_));
 sky130_fd_sc_hd__nand3_4 _34649_ (.A(_06357_),
    .B(_06895_),
    .C(_20107_),
    .Y(_12087_));
 sky130_fd_sc_hd__nor2_8 _34650_ (.A(_08037_),
    .B(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a22o_2 _34651_ (.A1(_11486_),
    .A2(_08453_),
    .B1(_07115_),
    .B2(_08884_),
    .X(_12089_));
 sky130_fd_sc_hd__nand2_4 _34652_ (.A(net505),
    .B(_20101_),
    .Y(_12090_));
 sky130_vsdinv _34653_ (.A(_12090_),
    .Y(_12091_));
 sky130_fd_sc_hd__nand2_1 _34654_ (.A(_12089_),
    .B(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__buf_6 _34655_ (.A(_11734_),
    .X(_12093_));
 sky130_fd_sc_hd__o22ai_4 _34656_ (.A1(_12093_),
    .A2(_11721_),
    .B1(_11725_),
    .B2(_11728_),
    .Y(_12094_));
 sky130_fd_sc_hd__a22oi_4 _34657_ (.A1(net444),
    .A2(_20108_),
    .B1(_10351_),
    .B2(_11078_),
    .Y(_12095_));
 sky130_fd_sc_hd__o21ai_2 _34658_ (.A1(_12095_),
    .A2(_12088_),
    .B1(_12090_),
    .Y(_12096_));
 sky130_fd_sc_hd__o211ai_4 _34659_ (.A1(_12088_),
    .A2(_12092_),
    .B1(_12094_),
    .C1(_12096_),
    .Y(_12097_));
 sky130_fd_sc_hd__o21ai_4 _34660_ (.A1(_12095_),
    .A2(_12088_),
    .B1(_12091_),
    .Y(_12098_));
 sky130_fd_sc_hd__o22a_4 _34661_ (.A1(_09733_),
    .A2(_11721_),
    .B1(_11725_),
    .B2(_11728_),
    .X(_12099_));
 sky130_fd_sc_hd__buf_6 _34662_ (.A(_08037_),
    .X(_12100_));
 sky130_fd_sc_hd__o211ai_4 _34663_ (.A1(_12100_),
    .A2(_12087_),
    .B1(_12090_),
    .C1(_12089_),
    .Y(_12101_));
 sky130_fd_sc_hd__buf_4 _34664_ (.A(_09037_),
    .X(_12102_));
 sky130_fd_sc_hd__buf_4 _34665_ (.A(_20096_),
    .X(_12103_));
 sky130_fd_sc_hd__nand2_8 _34666_ (.A(_12102_),
    .B(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__nor2_8 _34667_ (.A(_06623_),
    .B(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__nand2_2 _34668_ (.A(_05953_),
    .B(_09487_),
    .Y(_12106_));
 sky130_fd_sc_hd__a22o_2 _34669_ (.A1(_10337_),
    .A2(_11205_),
    .B1(_06046_),
    .B2(_20094_),
    .X(_12107_));
 sky130_fd_sc_hd__nand3b_4 _34670_ (.A_N(_12105_),
    .B(_12106_),
    .C(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__buf_4 _34671_ (.A(_09038_),
    .X(_12109_));
 sky130_fd_sc_hd__a22oi_4 _34672_ (.A1(_06119_),
    .A2(_11205_),
    .B1(_06046_),
    .B2(_12109_),
    .Y(_12110_));
 sky130_vsdinv _34673_ (.A(_12106_),
    .Y(_12111_));
 sky130_fd_sc_hd__o21ai_2 _34674_ (.A1(_12110_),
    .A2(_12105_),
    .B1(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__a32oi_4 _34675_ (.A1(_12098_),
    .A2(_12099_),
    .A3(_12101_),
    .B1(_12108_),
    .B2(_12112_),
    .Y(_12113_));
 sky130_fd_sc_hd__nand3_4 _34676_ (.A(_12098_),
    .B(_12099_),
    .C(_12101_),
    .Y(_12114_));
 sky130_fd_sc_hd__nand2_2 _34677_ (.A(_12108_),
    .B(_12112_),
    .Y(_12115_));
 sky130_fd_sc_hd__a21oi_4 _34678_ (.A1(_12097_),
    .A2(_12114_),
    .B1(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__a21oi_4 _34679_ (.A1(_12097_),
    .A2(_12113_),
    .B1(_12116_),
    .Y(_12117_));
 sky130_fd_sc_hd__a21oi_2 _34680_ (.A1(_12081_),
    .A2(_12086_),
    .B1(_12117_),
    .Y(_12118_));
 sky130_fd_sc_hd__o2bb2ai_1 _34681_ (.A1_N(_12084_),
    .A2_N(_12083_),
    .B1(_11708_),
    .B2(_11712_),
    .Y(_12119_));
 sky130_fd_sc_hd__o211a_1 _34682_ (.A1(_12080_),
    .A2(_12119_),
    .B1(_12117_),
    .C1(_12081_),
    .X(_12120_));
 sky130_fd_sc_hd__o22ai_4 _34683_ (.A1(_11892_),
    .A2(_12057_),
    .B1(_12118_),
    .B2(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__o21ai_4 _34684_ (.A1(_11895_),
    .A2(_11892_),
    .B1(_11887_),
    .Y(_12122_));
 sky130_fd_sc_hd__a21oi_4 _34685_ (.A1(_12098_),
    .A2(_12101_),
    .B1(_12099_),
    .Y(_12123_));
 sky130_fd_sc_hd__nand2_2 _34686_ (.A(_12114_),
    .B(_12115_),
    .Y(_12124_));
 sky130_fd_sc_hd__nor2_4 _34687_ (.A(_12123_),
    .B(_12124_),
    .Y(_12125_));
 sky130_fd_sc_hd__o2bb2ai_4 _34688_ (.A1_N(_12086_),
    .A2_N(_12081_),
    .B1(_12116_),
    .B2(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__nand3_4 _34689_ (.A(_12081_),
    .B(_12086_),
    .C(_12117_),
    .Y(_12127_));
 sky130_fd_sc_hd__nand3_4 _34690_ (.A(_12122_),
    .B(_12126_),
    .C(_12127_),
    .Y(_12128_));
 sky130_fd_sc_hd__nand2_1 _34691_ (.A(_11755_),
    .B(_11720_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand2_4 _34692_ (.A(_12129_),
    .B(_11717_),
    .Y(_12130_));
 sky130_fd_sc_hd__nand3_2 _34693_ (.A(_12121_),
    .B(_12128_),
    .C(_12130_),
    .Y(_12131_));
 sky130_vsdinv _34694_ (.A(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__a21oi_4 _34695_ (.A1(_12121_),
    .A2(_12128_),
    .B1(_12130_),
    .Y(_12133_));
 sky130_fd_sc_hd__nand2_2 _34696_ (.A(_11813_),
    .B(_11844_),
    .Y(_12134_));
 sky130_fd_sc_hd__nand2_1 _34697_ (.A(_12134_),
    .B(_11820_),
    .Y(_12135_));
 sky130_fd_sc_hd__nand3_4 _34698_ (.A(_10961_),
    .B(_10962_),
    .C(_20164_),
    .Y(_12136_));
 sky130_fd_sc_hd__nor2_2 _34699_ (.A(_06614_),
    .B(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__a22oi_4 _34700_ (.A1(_11777_),
    .A2(_05244_),
    .B1(_05369_),
    .B2(_18693_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand2_4 _34701_ (.A(_19832_),
    .B(_05285_),
    .Y(_12139_));
 sky130_vsdinv _34702_ (.A(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__o21ai_2 _34703_ (.A1(_12137_),
    .A2(_12138_),
    .B1(_12140_),
    .Y(_12141_));
 sky130_fd_sc_hd__o2bb2ai_4 _34704_ (.A1_N(_11777_),
    .A2_N(_06199_),
    .B1(_05182_),
    .B2(_10967_),
    .Y(_12142_));
 sky130_fd_sc_hd__o211ai_4 _34705_ (.A1(_20169_),
    .A2(_12136_),
    .B1(_12139_),
    .C1(_12142_),
    .Y(_12143_));
 sky130_fd_sc_hd__o21ai_1 _34706_ (.A1(_06197_),
    .A2(_11775_),
    .B1(_11780_),
    .Y(_12144_));
 sky130_fd_sc_hd__nand2_2 _34707_ (.A(_12144_),
    .B(_11784_),
    .Y(_12145_));
 sky130_fd_sc_hd__nand3_4 _34708_ (.A(_12141_),
    .B(_12143_),
    .C(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__o21ai_2 _34709_ (.A1(_12137_),
    .A2(_12138_),
    .B1(_12139_),
    .Y(_12147_));
 sky130_fd_sc_hd__o211ai_4 _34710_ (.A1(_05183_),
    .A2(_12136_),
    .B1(_12140_),
    .C1(_12142_),
    .Y(_12148_));
 sky130_fd_sc_hd__o22ai_4 _34711_ (.A1(_05144_),
    .A2(_11775_),
    .B1(_11780_),
    .B2(_11779_),
    .Y(_12149_));
 sky130_fd_sc_hd__nand3_4 _34712_ (.A(_12147_),
    .B(_12148_),
    .C(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__nand2_1 _34713_ (.A(_12146_),
    .B(_12150_),
    .Y(_12151_));
 sky130_fd_sc_hd__nand2_4 _34714_ (.A(_05696_),
    .B(_05391_),
    .Y(_12152_));
 sky130_fd_sc_hd__nor2_8 _34715_ (.A(_10983_),
    .B(_12152_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_2 _34716_ (.A(_09696_),
    .B(_05698_),
    .Y(_12154_));
 sky130_fd_sc_hd__a22o_2 _34717_ (.A1(_10411_),
    .A2(_05577_),
    .B1(_10412_),
    .B2(_05693_),
    .X(_12155_));
 sky130_fd_sc_hd__nand3b_2 _34718_ (.A_N(_12153_),
    .B(_12154_),
    .C(_12155_),
    .Y(_12156_));
 sky130_fd_sc_hd__a22oi_4 _34719_ (.A1(_09997_),
    .A2(_05577_),
    .B1(_09998_),
    .B2(_05697_),
    .Y(_12157_));
 sky130_vsdinv _34720_ (.A(_12154_),
    .Y(_12158_));
 sky130_fd_sc_hd__o21ai_2 _34721_ (.A1(_12157_),
    .A2(_12153_),
    .B1(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__nand2_4 _34722_ (.A(_12156_),
    .B(_12159_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand2_2 _34723_ (.A(_12151_),
    .B(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__a21boi_2 _34724_ (.A1(_11788_),
    .A2(_11817_),
    .B1_N(_11792_),
    .Y(_12162_));
 sky130_fd_sc_hd__nand2_1 _34725_ (.A(_12155_),
    .B(_12158_),
    .Y(_12163_));
 sky130_fd_sc_hd__o21ai_1 _34726_ (.A1(_12157_),
    .A2(_12153_),
    .B1(_12154_),
    .Y(_12164_));
 sky130_fd_sc_hd__o21ai_2 _34727_ (.A1(_12153_),
    .A2(_12163_),
    .B1(_12164_),
    .Y(_12165_));
 sky130_fd_sc_hd__nand3_4 _34728_ (.A(_12146_),
    .B(_12150_),
    .C(_12165_),
    .Y(_12166_));
 sky130_fd_sc_hd__nand3_4 _34729_ (.A(_12161_),
    .B(_12162_),
    .C(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__nand2_1 _34730_ (.A(_12151_),
    .B(_12165_),
    .Y(_12168_));
 sky130_fd_sc_hd__nand2_2 _34731_ (.A(_11788_),
    .B(_11817_),
    .Y(_12169_));
 sky130_fd_sc_hd__nand2_1 _34732_ (.A(_12169_),
    .B(_11793_),
    .Y(_12170_));
 sky130_fd_sc_hd__nand3_2 _34733_ (.A(_12146_),
    .B(_12150_),
    .C(_12160_),
    .Y(_12171_));
 sky130_fd_sc_hd__nand3_4 _34734_ (.A(_12168_),
    .B(_12170_),
    .C(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__a22oi_4 _34735_ (.A1(_10552_),
    .A2(_05820_),
    .B1(_11010_),
    .B2(_05823_),
    .Y(_12173_));
 sky130_fd_sc_hd__nand3_4 _34736_ (.A(_11008_),
    .B(_09981_),
    .C(_05699_),
    .Y(_12174_));
 sky130_fd_sc_hd__nor2_8 _34737_ (.A(net445),
    .B(_12174_),
    .Y(_12175_));
 sky130_fd_sc_hd__nand2_2 _34738_ (.A(_19853_),
    .B(_07024_),
    .Y(_12176_));
 sky130_vsdinv _34739_ (.A(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__o21ai_4 _34740_ (.A1(_12173_),
    .A2(_12175_),
    .B1(_12177_),
    .Y(_12178_));
 sky130_fd_sc_hd__a21oi_4 _34741_ (.A1(_11802_),
    .A2(_11798_),
    .B1(_11796_),
    .Y(_12179_));
 sky130_fd_sc_hd__a22o_2 _34742_ (.A1(_11826_),
    .A2(_06289_),
    .B1(_10384_),
    .B2(_20146_),
    .X(_12180_));
 sky130_fd_sc_hd__o211ai_4 _34743_ (.A1(_06288_),
    .A2(_12174_),
    .B1(_12176_),
    .C1(_12180_),
    .Y(_12181_));
 sky130_fd_sc_hd__nand3_4 _34744_ (.A(_12178_),
    .B(_12179_),
    .C(_12181_),
    .Y(_12182_));
 sky130_fd_sc_hd__o21ai_2 _34745_ (.A1(_12173_),
    .A2(_12175_),
    .B1(_12176_),
    .Y(_12183_));
 sky130_fd_sc_hd__o211ai_4 _34746_ (.A1(_06288_),
    .A2(_12174_),
    .B1(_12177_),
    .C1(_12180_),
    .Y(_12184_));
 sky130_fd_sc_hd__o22ai_4 _34747_ (.A1(_06624_),
    .A2(net440),
    .B1(_11797_),
    .B2(_11795_),
    .Y(_12185_));
 sky130_fd_sc_hd__nand3_4 _34748_ (.A(_12183_),
    .B(_12184_),
    .C(_12185_),
    .Y(_12186_));
 sky130_fd_sc_hd__o21ai_4 _34749_ (.A1(_11823_),
    .A2(_11821_),
    .B1(_11830_),
    .Y(_12187_));
 sky130_fd_sc_hd__and3_1 _34750_ (.A(_12182_),
    .B(_12186_),
    .C(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__a21oi_4 _34751_ (.A1(_12182_),
    .A2(_12186_),
    .B1(_12187_),
    .Y(_12189_));
 sky130_fd_sc_hd__o2bb2ai_2 _34752_ (.A1_N(_12167_),
    .A2_N(_12172_),
    .B1(_12188_),
    .B2(_12189_),
    .Y(_12190_));
 sky130_fd_sc_hd__o21a_1 _34753_ (.A1(_11823_),
    .A2(_11821_),
    .B1(_11830_),
    .X(_12191_));
 sky130_fd_sc_hd__a31oi_4 _34754_ (.A1(_12179_),
    .A2(_12178_),
    .A3(_12181_),
    .B1(_12191_),
    .Y(_12192_));
 sky130_fd_sc_hd__a21oi_4 _34755_ (.A1(_12186_),
    .A2(_12192_),
    .B1(_12189_),
    .Y(_12193_));
 sky130_fd_sc_hd__nand3_4 _34756_ (.A(_12172_),
    .B(_12167_),
    .C(_12193_),
    .Y(_12194_));
 sky130_fd_sc_hd__nand3_4 _34757_ (.A(_12135_),
    .B(_12190_),
    .C(_12194_),
    .Y(_12195_));
 sky130_fd_sc_hd__nand2_2 _34758_ (.A(_12172_),
    .B(_12167_),
    .Y(_12196_));
 sky130_fd_sc_hd__nand2_4 _34759_ (.A(_12196_),
    .B(_12193_),
    .Y(_12197_));
 sky130_fd_sc_hd__a21boi_4 _34760_ (.A1(_11813_),
    .A2(_11844_),
    .B1_N(_11819_),
    .Y(_12198_));
 sky130_fd_sc_hd__a21o_2 _34761_ (.A1(_12186_),
    .A2(_12192_),
    .B1(_12189_),
    .X(_12199_));
 sky130_fd_sc_hd__nand3_4 _34762_ (.A(_12199_),
    .B(_12172_),
    .C(_12167_),
    .Y(_12200_));
 sky130_fd_sc_hd__nand3_4 _34763_ (.A(_12197_),
    .B(_12198_),
    .C(_12200_),
    .Y(_12201_));
 sky130_fd_sc_hd__a22oi_4 _34764_ (.A1(_10916_),
    .A2(_05986_),
    .B1(_07965_),
    .B2(_06143_),
    .Y(_12202_));
 sky130_fd_sc_hd__and4_2 _34765_ (.A(_08582_),
    .B(_08577_),
    .C(_06438_),
    .D(_07502_),
    .X(_12203_));
 sky130_fd_sc_hd__nand2_4 _34766_ (.A(_19865_),
    .B(_06989_),
    .Y(_12204_));
 sky130_vsdinv _34767_ (.A(_12204_),
    .Y(_12205_));
 sky130_fd_sc_hd__o21ai_2 _34768_ (.A1(_12202_),
    .A2(_12203_),
    .B1(_12205_),
    .Y(_12206_));
 sky130_fd_sc_hd__a21oi_2 _34769_ (.A1(_11854_),
    .A2(_11856_),
    .B1(_11853_),
    .Y(_12207_));
 sky130_fd_sc_hd__nand2_1 _34770_ (.A(_19858_),
    .B(_06696_),
    .Y(_12208_));
 sky130_fd_sc_hd__nand3b_4 _34771_ (.A_N(_12208_),
    .B(_08592_),
    .C(_07004_),
    .Y(_12209_));
 sky130_fd_sc_hd__a22o_1 _34772_ (.A1(_10916_),
    .A2(_05986_),
    .B1(_08775_),
    .B2(_06442_),
    .X(_12210_));
 sky130_fd_sc_hd__nand3_2 _34773_ (.A(_12209_),
    .B(_12210_),
    .C(_12204_),
    .Y(_12211_));
 sky130_fd_sc_hd__nand3_4 _34774_ (.A(_12206_),
    .B(_12207_),
    .C(_12211_),
    .Y(_12212_));
 sky130_fd_sc_hd__o21ai_2 _34775_ (.A1(_12202_),
    .A2(_12203_),
    .B1(_12204_),
    .Y(_12213_));
 sky130_fd_sc_hd__nand3_2 _34776_ (.A(_12209_),
    .B(_12210_),
    .C(_12205_),
    .Y(_12214_));
 sky130_fd_sc_hd__o22ai_4 _34777_ (.A1(net465),
    .A2(_11852_),
    .B1(_11855_),
    .B2(_11859_),
    .Y(_12215_));
 sky130_fd_sc_hd__nand3_4 _34778_ (.A(_12213_),
    .B(_12214_),
    .C(_12215_),
    .Y(_12216_));
 sky130_fd_sc_hd__nand2_1 _34779_ (.A(_12212_),
    .B(_12216_),
    .Y(_12217_));
 sky130_fd_sc_hd__a22oi_4 _34780_ (.A1(_08779_),
    .A2(_20129_),
    .B1(_08598_),
    .B2(_07257_),
    .Y(_12218_));
 sky130_fd_sc_hd__nand2_8 _34781_ (.A(_08326_),
    .B(_19873_),
    .Y(_12219_));
 sky130_fd_sc_hd__nor2_4 _34782_ (.A(_08144_),
    .B(_12219_),
    .Y(_12220_));
 sky130_fd_sc_hd__nor2_1 _34783_ (.A(_12218_),
    .B(_12220_),
    .Y(_12221_));
 sky130_fd_sc_hd__nand2_4 _34784_ (.A(_07356_),
    .B(_07251_),
    .Y(_12222_));
 sky130_vsdinv _34785_ (.A(_12222_),
    .Y(_12223_));
 sky130_fd_sc_hd__nand2_1 _34786_ (.A(_12221_),
    .B(_12223_),
    .Y(_12224_));
 sky130_fd_sc_hd__o21ai_1 _34787_ (.A1(_12218_),
    .A2(_12220_),
    .B1(_12222_),
    .Y(_12225_));
 sky130_fd_sc_hd__nand2_1 _34788_ (.A(_12224_),
    .B(_12225_),
    .Y(_12226_));
 sky130_fd_sc_hd__nand2_1 _34789_ (.A(_12217_),
    .B(_12226_),
    .Y(_12227_));
 sky130_fd_sc_hd__nand2_1 _34790_ (.A(_12221_),
    .B(_12222_),
    .Y(_12228_));
 sky130_fd_sc_hd__o21ai_1 _34791_ (.A1(_12218_),
    .A2(_12220_),
    .B1(_12223_),
    .Y(_12229_));
 sky130_fd_sc_hd__nand2_1 _34792_ (.A(_12228_),
    .B(_12229_),
    .Y(_12230_));
 sky130_fd_sc_hd__nand3_4 _34793_ (.A(_12230_),
    .B(_12212_),
    .C(_12216_),
    .Y(_12231_));
 sky130_fd_sc_hd__o21ai_2 _34794_ (.A1(_11838_),
    .A2(_11839_),
    .B1(_11835_),
    .Y(_12232_));
 sky130_fd_sc_hd__nand3_4 _34795_ (.A(_12227_),
    .B(_12231_),
    .C(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__buf_2 _34796_ (.A(_12233_),
    .X(_12234_));
 sky130_vsdinv _34797_ (.A(_12229_),
    .Y(_12235_));
 sky130_fd_sc_hd__and2_1 _34798_ (.A(_12221_),
    .B(_12222_),
    .X(_12236_));
 sky130_fd_sc_hd__o2bb2ai_1 _34799_ (.A1_N(_12216_),
    .A2_N(_12212_),
    .B1(_12235_),
    .B2(_12236_),
    .Y(_12237_));
 sky130_fd_sc_hd__o21a_1 _34800_ (.A1(_11345_),
    .A2(_11356_),
    .B1(_11830_),
    .X(_12238_));
 sky130_fd_sc_hd__a22oi_2 _34801_ (.A1(_12238_),
    .A2(_11825_),
    .B1(_11833_),
    .B2(_11836_),
    .Y(_12239_));
 sky130_fd_sc_hd__nand3_1 _34802_ (.A(_12226_),
    .B(_12212_),
    .C(_12216_),
    .Y(_12240_));
 sky130_fd_sc_hd__nand3_2 _34803_ (.A(_12237_),
    .B(_12239_),
    .C(_12240_),
    .Y(_12241_));
 sky130_fd_sc_hd__clkbuf_4 _34804_ (.A(_12241_),
    .X(_12242_));
 sky130_vsdinv _34805_ (.A(_11865_),
    .Y(_12243_));
 sky130_fd_sc_hd__o21ai_4 _34806_ (.A1(_11879_),
    .A2(_12243_),
    .B1(_11861_),
    .Y(_12244_));
 sky130_fd_sc_hd__a21oi_4 _34807_ (.A1(_12234_),
    .A2(_12242_),
    .B1(_12244_),
    .Y(_12245_));
 sky130_fd_sc_hd__and3_4 _34808_ (.A(_12233_),
    .B(_12241_),
    .C(_12244_),
    .X(_12246_));
 sky130_fd_sc_hd__o2bb2ai_4 _34809_ (.A1_N(_12195_),
    .A2_N(_12201_),
    .B1(_12245_),
    .B2(_12246_),
    .Y(_12247_));
 sky130_fd_sc_hd__nor2_8 _34810_ (.A(_12245_),
    .B(_12246_),
    .Y(_12248_));
 sky130_fd_sc_hd__nand3_4 _34811_ (.A(_12201_),
    .B(_12195_),
    .C(_12248_),
    .Y(_12249_));
 sky130_vsdinv _34812_ (.A(_11845_),
    .Y(_12250_));
 sky130_fd_sc_hd__nand2_1 _34813_ (.A(_11774_),
    .B(_11843_),
    .Y(_12251_));
 sky130_fd_sc_hd__o2bb2ai_4 _34814_ (.A1_N(_11851_),
    .A2_N(_11897_),
    .B1(_12250_),
    .B2(_12251_),
    .Y(_12252_));
 sky130_fd_sc_hd__a21oi_4 _34815_ (.A1(_12247_),
    .A2(_12249_),
    .B1(_12252_),
    .Y(_12253_));
 sky130_fd_sc_hd__a21oi_4 _34816_ (.A1(_12197_),
    .A2(_12200_),
    .B1(_12198_),
    .Y(_12254_));
 sky130_fd_sc_hd__nand2_1 _34817_ (.A(_12201_),
    .B(_12248_),
    .Y(_12255_));
 sky130_fd_sc_hd__o211a_2 _34818_ (.A1(_12254_),
    .A2(_12255_),
    .B1(_12247_),
    .C1(_12252_),
    .X(_12256_));
 sky130_fd_sc_hd__o22ai_4 _34819_ (.A1(_12132_),
    .A2(_12133_),
    .B1(_12253_),
    .B2(_12256_),
    .Y(_12257_));
 sky130_fd_sc_hd__a2bb2oi_2 _34820_ (.A1_N(_12245_),
    .A2_N(_12246_),
    .B1(_12195_),
    .B2(_12201_),
    .Y(_12258_));
 sky130_vsdinv _34821_ (.A(_11861_),
    .Y(_12259_));
 sky130_fd_sc_hd__a21oi_1 _34822_ (.A1(_11883_),
    .A2(_11865_),
    .B1(_12259_),
    .Y(_12260_));
 sky130_fd_sc_hd__and3_1 _34823_ (.A(_12234_),
    .B(_12242_),
    .C(_12260_),
    .X(_12261_));
 sky130_fd_sc_hd__a21oi_1 _34824_ (.A1(_12234_),
    .A2(_12242_),
    .B1(_12260_),
    .Y(_12262_));
 sky130_fd_sc_hd__o211a_4 _34825_ (.A1(_12261_),
    .A2(_12262_),
    .B1(_12195_),
    .C1(_12201_),
    .X(_12263_));
 sky130_fd_sc_hd__a21boi_2 _34826_ (.A1(_11897_),
    .A2(_11851_),
    .B1_N(_11846_),
    .Y(_12264_));
 sky130_fd_sc_hd__o21ai_4 _34827_ (.A1(_12258_),
    .A2(_12263_),
    .B1(_12264_),
    .Y(_12265_));
 sky130_fd_sc_hd__nand2_1 _34828_ (.A(_12126_),
    .B(_12127_),
    .Y(_12266_));
 sky130_fd_sc_hd__a21oi_4 _34829_ (.A1(_11886_),
    .A2(_11888_),
    .B1(_11893_),
    .Y(_12267_));
 sky130_fd_sc_hd__a21boi_4 _34830_ (.A1(_12266_),
    .A2(_12267_),
    .B1_N(_12130_),
    .Y(_12268_));
 sky130_fd_sc_hd__a21oi_4 _34831_ (.A1(_12128_),
    .A2(_12268_),
    .B1(_12133_),
    .Y(_12269_));
 sky130_fd_sc_hd__nand3_4 _34832_ (.A(_12252_),
    .B(_12247_),
    .C(_12249_),
    .Y(_12270_));
 sky130_fd_sc_hd__nand3_4 _34833_ (.A(_12265_),
    .B(_12269_),
    .C(_12270_),
    .Y(_12271_));
 sky130_fd_sc_hd__o21ai_4 _34834_ (.A1(_11924_),
    .A2(_11901_),
    .B1(_11913_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand3_4 _34835_ (.A(_12257_),
    .B(_12271_),
    .C(_12272_),
    .Y(_12273_));
 sky130_fd_sc_hd__o21ai_2 _34836_ (.A1(_12253_),
    .A2(_12256_),
    .B1(_12269_),
    .Y(_12274_));
 sky130_fd_sc_hd__a21oi_4 _34837_ (.A1(_11912_),
    .A2(_11915_),
    .B1(_11905_),
    .Y(_12275_));
 sky130_fd_sc_hd__a21oi_4 _34838_ (.A1(_12126_),
    .A2(_12127_),
    .B1(_12122_),
    .Y(_12276_));
 sky130_vsdinv _34839_ (.A(_12086_),
    .Y(_12277_));
 sky130_fd_sc_hd__nand2_2 _34840_ (.A(_12081_),
    .B(_12117_),
    .Y(_12278_));
 sky130_fd_sc_hd__o211a_1 _34841_ (.A1(_12277_),
    .A2(_12278_),
    .B1(_12126_),
    .C1(_12122_),
    .X(_12279_));
 sky130_vsdinv _34842_ (.A(_12130_),
    .Y(_12280_));
 sky130_fd_sc_hd__o21ai_1 _34843_ (.A1(_12276_),
    .A2(_12279_),
    .B1(_12280_),
    .Y(_12281_));
 sky130_fd_sc_hd__nand2_2 _34844_ (.A(_12281_),
    .B(_12131_),
    .Y(_12282_));
 sky130_fd_sc_hd__nand3_2 _34845_ (.A(_12265_),
    .B(_12270_),
    .C(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__nand3_4 _34846_ (.A(_12274_),
    .B(_12275_),
    .C(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__o21a_1 _34847_ (.A1(_11954_),
    .A2(_11949_),
    .B1(_11955_),
    .X(_12285_));
 sky130_vsdinv _34848_ (.A(_11938_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand2_1 _34849_ (.A(_11943_),
    .B(_11946_),
    .Y(_12287_));
 sky130_vsdinv _34850_ (.A(_12287_),
    .Y(_12288_));
 sky130_fd_sc_hd__nand2_2 _34851_ (.A(_11731_),
    .B(_11751_),
    .Y(_12289_));
 sky130_fd_sc_hd__a22oi_4 _34852_ (.A1(_19913_),
    .A2(_11934_),
    .B1(_19916_),
    .B2(_11157_),
    .Y(_12290_));
 sky130_fd_sc_hd__nand3_4 _34853_ (.A(_06483_),
    .B(_06657_),
    .C(_10259_),
    .Y(_12291_));
 sky130_fd_sc_hd__nor2_8 _34854_ (.A(_10265_),
    .B(_12291_),
    .Y(_12292_));
 sky130_fd_sc_hd__nand2_2 _34855_ (.A(_19918_),
    .B(_20078_),
    .Y(_12293_));
 sky130_vsdinv _34856_ (.A(_12293_),
    .Y(_12294_));
 sky130_fd_sc_hd__o21ai_2 _34857_ (.A1(_12290_),
    .A2(_12292_),
    .B1(_12294_),
    .Y(_12295_));
 sky130_fd_sc_hd__a21oi_2 _34858_ (.A1(_11738_),
    .A2(_11741_),
    .B1(_11743_),
    .Y(_12296_));
 sky130_fd_sc_hd__buf_6 _34859_ (.A(_10265_),
    .X(_12297_));
 sky130_fd_sc_hd__buf_4 _34860_ (.A(_10259_),
    .X(_12298_));
 sky130_fd_sc_hd__a22o_2 _34861_ (.A1(_19913_),
    .A2(_10262_),
    .B1(_19916_),
    .B2(_12298_),
    .X(_12299_));
 sky130_fd_sc_hd__o211ai_4 _34862_ (.A1(_12297_),
    .A2(_12291_),
    .B1(_12293_),
    .C1(_12299_),
    .Y(_12300_));
 sky130_fd_sc_hd__nand3_4 _34863_ (.A(_12295_),
    .B(_12296_),
    .C(_12300_),
    .Y(_12301_));
 sky130_fd_sc_hd__o21ai_2 _34864_ (.A1(_12290_),
    .A2(_12292_),
    .B1(_12293_),
    .Y(_12302_));
 sky130_fd_sc_hd__buf_4 _34865_ (.A(_08881_),
    .X(_12303_));
 sky130_fd_sc_hd__buf_4 _34866_ (.A(_11503_),
    .X(_12304_));
 sky130_fd_sc_hd__a22oi_4 _34867_ (.A1(_19903_),
    .A2(_12303_),
    .B1(_19907_),
    .B2(_12304_),
    .Y(_12305_));
 sky130_fd_sc_hd__o22ai_4 _34868_ (.A1(_06623_),
    .A2(_11737_),
    .B1(_11740_),
    .B2(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__buf_6 _34869_ (.A(_10265_),
    .X(_12307_));
 sky130_fd_sc_hd__o211ai_2 _34870_ (.A1(_12307_),
    .A2(_12291_),
    .B1(_12294_),
    .C1(_12299_),
    .Y(_12308_));
 sky130_fd_sc_hd__nand3_4 _34871_ (.A(_12302_),
    .B(_12306_),
    .C(_12308_),
    .Y(_12309_));
 sky130_fd_sc_hd__a21o_2 _34872_ (.A1(_11935_),
    .A2(_11933_),
    .B1(_11930_),
    .X(_12310_));
 sky130_fd_sc_hd__a21o_2 _34873_ (.A1(_12301_),
    .A2(_12309_),
    .B1(_12310_),
    .X(_12311_));
 sky130_fd_sc_hd__nand3_4 _34874_ (.A(_12301_),
    .B(_12309_),
    .C(_12310_),
    .Y(_12312_));
 sky130_fd_sc_hd__a22oi_4 _34875_ (.A1(_11736_),
    .A2(_12289_),
    .B1(_12311_),
    .B2(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__a21oi_4 _34876_ (.A1(_11732_),
    .A2(_11735_),
    .B1(_11733_),
    .Y(_12314_));
 sky130_fd_sc_hd__a32oi_4 _34877_ (.A1(_11732_),
    .A2(_11733_),
    .A3(_11735_),
    .B1(_11742_),
    .B2(_11744_),
    .Y(_12315_));
 sky130_fd_sc_hd__o211a_2 _34878_ (.A1(_12314_),
    .A2(_12315_),
    .B1(_12312_),
    .C1(_12311_),
    .X(_12316_));
 sky130_fd_sc_hd__o22ai_4 _34879_ (.A1(_12286_),
    .A2(_12288_),
    .B1(_12313_),
    .B2(_12316_),
    .Y(_12317_));
 sky130_fd_sc_hd__a22o_2 _34880_ (.A1(_11736_),
    .A2(_12289_),
    .B1(_12311_),
    .B2(_12312_),
    .X(_12318_));
 sky130_fd_sc_hd__o211ai_4 _34881_ (.A1(_12314_),
    .A2(_12315_),
    .B1(_12312_),
    .C1(_12311_),
    .Y(_12319_));
 sky130_fd_sc_hd__nand2_1 _34882_ (.A(_12287_),
    .B(_11938_),
    .Y(_12320_));
 sky130_vsdinv _34883_ (.A(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__nand3_2 _34884_ (.A(_12318_),
    .B(_12319_),
    .C(_12321_),
    .Y(_12322_));
 sky130_fd_sc_hd__nand3_4 _34885_ (.A(_12285_),
    .B(_12317_),
    .C(_12322_),
    .Y(_12323_));
 sky130_vsdinv _34886_ (.A(_11943_),
    .Y(_12324_));
 sky130_fd_sc_hd__nor2_2 _34887_ (.A(_11946_),
    .B(_12286_),
    .Y(_12325_));
 sky130_fd_sc_hd__o22ai_4 _34888_ (.A1(_12324_),
    .A2(_12325_),
    .B1(_12313_),
    .B2(_12316_),
    .Y(_12326_));
 sky130_fd_sc_hd__nand3_2 _34889_ (.A(_12318_),
    .B(_12319_),
    .C(_12320_),
    .Y(_12327_));
 sky130_fd_sc_hd__o21ai_2 _34890_ (.A1(_11954_),
    .A2(_11949_),
    .B1(_11955_),
    .Y(_12328_));
 sky130_fd_sc_hd__nand3_4 _34891_ (.A(_12326_),
    .B(_12327_),
    .C(_12328_),
    .Y(_12329_));
 sky130_vsdinv _34892_ (.A(_11976_),
    .Y(_12330_));
 sky130_fd_sc_hd__and3_1 _34893_ (.A(_11974_),
    .B(_19929_),
    .C(_20071_),
    .X(_12331_));
 sky130_fd_sc_hd__nand2_1 _34894_ (.A(_11978_),
    .B(_11968_),
    .Y(_12332_));
 sky130_fd_sc_hd__nand2_1 _34895_ (.A(_12332_),
    .B(_11972_),
    .Y(_12333_));
 sky130_fd_sc_hd__nor2_2 _34896_ (.A(_11160_),
    .B(_11962_),
    .Y(_12334_));
 sky130_fd_sc_hd__nand2_4 _34897_ (.A(_05213_),
    .B(_20072_),
    .Y(_12335_));
 sky130_fd_sc_hd__nand2_4 _34898_ (.A(_05558_),
    .B(\pcpi_mul.rs1[31] ),
    .Y(_12336_));
 sky130_fd_sc_hd__nor2_8 _34899_ (.A(_12335_),
    .B(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__nand2_2 _34900_ (.A(_12335_),
    .B(_12336_),
    .Y(_12338_));
 sky130_fd_sc_hd__nand2_1 _34901_ (.A(_11161_),
    .B(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__and2_1 _34902_ (.A(_12335_),
    .B(_12336_),
    .X(_12340_));
 sky130_fd_sc_hd__o21ai_2 _34903_ (.A1(_12337_),
    .A2(_12340_),
    .B1(_11168_),
    .Y(_12341_));
 sky130_fd_sc_hd__o221ai_4 _34904_ (.A1(_11964_),
    .A2(_12334_),
    .B1(_12337_),
    .B2(_12339_),
    .C1(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__o21ai_2 _34905_ (.A1(_12337_),
    .A2(_12340_),
    .B1(_11161_),
    .Y(_12343_));
 sky130_fd_sc_hd__nand3b_2 _34906_ (.A_N(_12337_),
    .B(_11168_),
    .C(_12338_),
    .Y(_12344_));
 sky130_fd_sc_hd__a21oi_2 _34907_ (.A1(_11969_),
    .A2(_11161_),
    .B1(_11964_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand3_4 _34908_ (.A(_12343_),
    .B(_12344_),
    .C(_12345_),
    .Y(_12346_));
 sky130_fd_sc_hd__nand2_1 _34909_ (.A(_12342_),
    .B(_12346_),
    .Y(_12347_));
 sky130_fd_sc_hd__buf_1 _34910_ (.A(\pcpi_mul.rs1[32] ),
    .X(_12348_));
 sky130_fd_sc_hd__nand2_2 _34911_ (.A(net503),
    .B(_05247_),
    .Y(_12349_));
 sky130_vsdinv _34912_ (.A(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__nand2_2 _34913_ (.A(_11977_),
    .B(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__nand3_4 _34914_ (.A(_11974_),
    .B(_11976_),
    .C(_12349_),
    .Y(_12352_));
 sky130_fd_sc_hd__and2_1 _34915_ (.A(_12351_),
    .B(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__nand2_1 _34916_ (.A(_12347_),
    .B(_12353_),
    .Y(_12354_));
 sky130_fd_sc_hd__nand2_4 _34917_ (.A(_12351_),
    .B(_12352_),
    .Y(_12355_));
 sky130_fd_sc_hd__buf_2 _34918_ (.A(_12355_),
    .X(_12356_));
 sky130_fd_sc_hd__nand3_2 _34919_ (.A(_12342_),
    .B(_12346_),
    .C(_12356_),
    .Y(_12357_));
 sky130_fd_sc_hd__nand3_4 _34920_ (.A(_12333_),
    .B(_12354_),
    .C(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__o21a_1 _34921_ (.A1(_12330_),
    .A2(_12331_),
    .B1(_12358_),
    .X(_12359_));
 sky130_fd_sc_hd__a21boi_2 _34922_ (.A1(_11978_),
    .A2(_11968_),
    .B1_N(_11972_),
    .Y(_12360_));
 sky130_fd_sc_hd__nand2_1 _34923_ (.A(_12347_),
    .B(_12356_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand3_2 _34924_ (.A(_12342_),
    .B(_12353_),
    .C(_12346_),
    .Y(_12362_));
 sky130_fd_sc_hd__nand3_4 _34925_ (.A(_12360_),
    .B(_12361_),
    .C(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__nor2_1 _34926_ (.A(_12330_),
    .B(_12331_),
    .Y(_12364_));
 sky130_vsdinv _34927_ (.A(_12364_),
    .Y(_12365_));
 sky130_fd_sc_hd__a21oi_2 _34928_ (.A1(_12358_),
    .A2(_12363_),
    .B1(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__a21oi_4 _34929_ (.A1(_12359_),
    .A2(_12363_),
    .B1(_12366_),
    .Y(_12367_));
 sky130_fd_sc_hd__a21oi_4 _34930_ (.A1(_12323_),
    .A2(_12329_),
    .B1(_12367_),
    .Y(_12368_));
 sky130_vsdinv _34931_ (.A(_12363_),
    .Y(_12369_));
 sky130_fd_sc_hd__nand2_1 _34932_ (.A(_12358_),
    .B(_12365_),
    .Y(_12370_));
 sky130_fd_sc_hd__a21o_1 _34933_ (.A1(_12358_),
    .A2(_12363_),
    .B1(_12365_),
    .X(_12371_));
 sky130_fd_sc_hd__o2111a_1 _34934_ (.A1(_12369_),
    .A2(_12370_),
    .B1(_12371_),
    .C1(_12329_),
    .D1(_12323_),
    .X(_12372_));
 sky130_vsdinv _34935_ (.A(_11758_),
    .Y(_12373_));
 sky130_fd_sc_hd__nor2_4 _34936_ (.A(_12373_),
    .B(_11914_),
    .Y(_12374_));
 sky130_fd_sc_hd__o21ai_4 _34937_ (.A1(_12368_),
    .A2(_12372_),
    .B1(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__nand3_4 _34938_ (.A(_12367_),
    .B(_12323_),
    .C(_12329_),
    .Y(_12376_));
 sky130_fd_sc_hd__a21o_1 _34939_ (.A1(_12323_),
    .A2(_12329_),
    .B1(_12367_),
    .X(_12377_));
 sky130_fd_sc_hd__o211ai_4 _34940_ (.A1(_11914_),
    .A2(_12373_),
    .B1(_12376_),
    .C1(_12377_),
    .Y(_12378_));
 sky130_fd_sc_hd__a21bo_2 _34941_ (.A1(_11994_),
    .A2(_11957_),
    .B1_N(_11961_),
    .X(_12379_));
 sky130_fd_sc_hd__a21oi_4 _34942_ (.A1(_12375_),
    .A2(_12378_),
    .B1(_12379_),
    .Y(_12380_));
 sky130_fd_sc_hd__nand3_4 _34943_ (.A(_12375_),
    .B(_12378_),
    .C(_12379_),
    .Y(_12381_));
 sky130_vsdinv _34944_ (.A(_12381_),
    .Y(_12382_));
 sky130_fd_sc_hd__o2bb2ai_4 _34945_ (.A1_N(_12273_),
    .A2_N(_12284_),
    .B1(_12380_),
    .B2(_12382_),
    .Y(_12383_));
 sky130_fd_sc_hd__nand2_1 _34946_ (.A(_12377_),
    .B(_12376_),
    .Y(_12384_));
 sky130_fd_sc_hd__a21boi_4 _34947_ (.A1(_12384_),
    .A2(_12374_),
    .B1_N(_12379_),
    .Y(_12385_));
 sky130_fd_sc_hd__a21oi_4 _34948_ (.A1(_12378_),
    .A2(_12385_),
    .B1(_12380_),
    .Y(_12386_));
 sky130_fd_sc_hd__nand3_4 _34949_ (.A(_12386_),
    .B(_12273_),
    .C(_12284_),
    .Y(_12387_));
 sky130_fd_sc_hd__nand2_4 _34950_ (.A(_12025_),
    .B(_11919_),
    .Y(_12388_));
 sky130_fd_sc_hd__a21oi_4 _34951_ (.A1(_12383_),
    .A2(_12387_),
    .B1(_12388_),
    .Y(_12389_));
 sky130_fd_sc_hd__a32oi_2 _34952_ (.A1(_11920_),
    .A2(_11921_),
    .A3(_11925_),
    .B1(_12016_),
    .B2(_12018_),
    .Y(_12390_));
 sky130_fd_sc_hd__o211a_2 _34953_ (.A1(_12024_),
    .A2(_12390_),
    .B1(_12387_),
    .C1(_12383_),
    .X(_12391_));
 sky130_fd_sc_hd__nor2_4 _34954_ (.A(_11991_),
    .B(_12000_),
    .Y(_12392_));
 sky130_fd_sc_hd__a21oi_4 _34955_ (.A1(_12010_),
    .A2(_12005_),
    .B1(_12392_),
    .Y(_12393_));
 sky130_fd_sc_hd__and3_2 _34956_ (.A(_12010_),
    .B(_12005_),
    .C(_12392_),
    .X(_12394_));
 sky130_fd_sc_hd__nor2_8 _34957_ (.A(_12393_),
    .B(_12394_),
    .Y(_12395_));
 sky130_fd_sc_hd__o21ai_2 _34958_ (.A1(_12389_),
    .A2(_12391_),
    .B1(_12395_),
    .Y(_12396_));
 sky130_fd_sc_hd__nand2_1 _34959_ (.A(_11544_),
    .B(_11641_),
    .Y(_12397_));
 sky130_fd_sc_hd__a21oi_4 _34960_ (.A1(_11536_),
    .A2(_12397_),
    .B1(_12028_),
    .Y(_12398_));
 sky130_fd_sc_hd__a22oi_4 _34961_ (.A1(_12398_),
    .A2(_12020_),
    .B1(_12032_),
    .B2(_12041_),
    .Y(_12399_));
 sky130_fd_sc_hd__a21o_2 _34962_ (.A1(_12383_),
    .A2(_12387_),
    .B1(_12388_),
    .X(_12400_));
 sky130_vsdinv _34963_ (.A(_12395_),
    .Y(_12401_));
 sky130_fd_sc_hd__nand3_4 _34964_ (.A(_12388_),
    .B(_12387_),
    .C(_12383_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand3_2 _34965_ (.A(_12400_),
    .B(_12401_),
    .C(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__nand3_4 _34966_ (.A(_12396_),
    .B(_12399_),
    .C(_12403_),
    .Y(_12404_));
 sky130_fd_sc_hd__clkbuf_4 _34967_ (.A(_12393_),
    .X(_12405_));
 sky130_fd_sc_hd__o22ai_4 _34968_ (.A1(_12405_),
    .A2(_12394_),
    .B1(_12389_),
    .B2(_12391_),
    .Y(_12406_));
 sky130_fd_sc_hd__nand3_4 _34969_ (.A(_12400_),
    .B(_12395_),
    .C(_12402_),
    .Y(_12407_));
 sky130_fd_sc_hd__o21ai_2 _34970_ (.A1(_12034_),
    .A2(_12023_),
    .B1(_12033_),
    .Y(_12408_));
 sky130_fd_sc_hd__nand3_4 _34971_ (.A(_12406_),
    .B(_12407_),
    .C(_12408_),
    .Y(_12409_));
 sky130_fd_sc_hd__nand3_2 _34972_ (.A(_12404_),
    .B(_12409_),
    .C(_12037_),
    .Y(_12410_));
 sky130_vsdinv _34973_ (.A(_12410_),
    .Y(_12411_));
 sky130_vsdinv _34974_ (.A(_12037_),
    .Y(_12412_));
 sky130_fd_sc_hd__nand2_1 _34975_ (.A(_12404_),
    .B(_12409_),
    .Y(_12413_));
 sky130_fd_sc_hd__and3_1 _34976_ (.A(_12039_),
    .B(_12040_),
    .C(_12042_),
    .X(_12414_));
 sky130_vsdinv _34977_ (.A(_11668_),
    .Y(_12415_));
 sky130_fd_sc_hd__a31oi_2 _34978_ (.A1(_11686_),
    .A2(_12027_),
    .A3(_12035_),
    .B1(_12415_),
    .Y(_12416_));
 sky130_fd_sc_hd__o2bb2ai_2 _34979_ (.A1_N(_12412_),
    .A2_N(_12413_),
    .B1(_12414_),
    .B2(_12416_),
    .Y(_12417_));
 sky130_fd_sc_hd__o2bb2ai_1 _34980_ (.A1_N(_12409_),
    .A2_N(_12404_),
    .B1(_11688_),
    .B2(_11690_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand2_1 _34981_ (.A(_12036_),
    .B(_11668_),
    .Y(_12419_));
 sky130_fd_sc_hd__nand2_1 _34982_ (.A(_12419_),
    .B(_12043_),
    .Y(_12420_));
 sky130_fd_sc_hd__a21o_1 _34983_ (.A1(_12418_),
    .A2(_12410_),
    .B1(_12420_),
    .X(_12421_));
 sky130_fd_sc_hd__o21a_2 _34984_ (.A1(_12411_),
    .A2(_12417_),
    .B1(_12421_),
    .X(_12422_));
 sky130_fd_sc_hd__nand2_1 _34985_ (.A(_12056_),
    .B(_12051_),
    .Y(_12423_));
 sky130_fd_sc_hd__nand2_2 _34986_ (.A(_12423_),
    .B(_12048_),
    .Y(_12424_));
 sky130_fd_sc_hd__xnor2_4 _34987_ (.A(_12422_),
    .B(_12424_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21oi_4 _34988_ (.A1(_12400_),
    .A2(_12395_),
    .B1(_12391_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand2_1 _34989_ (.A(_12359_),
    .B(_12363_),
    .Y(_12426_));
 sky130_fd_sc_hd__nand2_4 _34990_ (.A(_12426_),
    .B(_12358_),
    .Y(_12427_));
 sky130_fd_sc_hd__nand2_2 _34991_ (.A(_12381_),
    .B(_12378_),
    .Y(_12428_));
 sky130_vsdinv _34992_ (.A(_12428_),
    .Y(_12429_));
 sky130_fd_sc_hd__nor2_4 _34993_ (.A(_12427_),
    .B(_12429_),
    .Y(_12430_));
 sky130_vsdinv _34994_ (.A(_12427_),
    .Y(_12431_));
 sky130_fd_sc_hd__nor2_4 _34995_ (.A(_12431_),
    .B(_12428_),
    .Y(_12432_));
 sky130_fd_sc_hd__nand2_2 _34996_ (.A(_12252_),
    .B(_12247_),
    .Y(_12433_));
 sky130_fd_sc_hd__o22ai_4 _34997_ (.A1(_12263_),
    .A2(_12433_),
    .B1(_12282_),
    .B2(_12253_),
    .Y(_12434_));
 sky130_fd_sc_hd__nor2_1 _34998_ (.A(_11883_),
    .B(_12259_),
    .Y(_12435_));
 sky130_fd_sc_hd__o2bb2ai_1 _34999_ (.A1_N(_12242_),
    .A2_N(_12234_),
    .B1(_12243_),
    .B2(_12435_),
    .Y(_12436_));
 sky130_fd_sc_hd__nand3_2 _35000_ (.A(_12233_),
    .B(_12242_),
    .C(_12244_),
    .Y(_12437_));
 sky130_fd_sc_hd__nand2_1 _35001_ (.A(_12436_),
    .B(_12437_),
    .Y(_12438_));
 sky130_fd_sc_hd__a31oi_4 _35002_ (.A1(_12197_),
    .A2(_12198_),
    .A3(_12200_),
    .B1(_12438_),
    .Y(_12439_));
 sky130_fd_sc_hd__a22oi_4 _35003_ (.A1(_10440_),
    .A2(_07004_),
    .B1(_19863_),
    .B2(_08546_),
    .Y(_12440_));
 sky130_fd_sc_hd__and4_2 _35004_ (.A(_10916_),
    .B(_08775_),
    .C(_20133_),
    .D(_20135_),
    .X(_12441_));
 sky130_fd_sc_hd__nand2_2 _35005_ (.A(_10435_),
    .B(_06813_),
    .Y(_12442_));
 sky130_vsdinv _35006_ (.A(_12442_),
    .Y(_12443_));
 sky130_fd_sc_hd__o21ai_2 _35007_ (.A1(_12440_),
    .A2(_12441_),
    .B1(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__a21oi_2 _35008_ (.A1(_12210_),
    .A2(_12205_),
    .B1(_12203_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand2_1 _35009_ (.A(_10916_),
    .B(_07503_),
    .Y(_12446_));
 sky130_fd_sc_hd__buf_6 _35010_ (.A(_08577_),
    .X(_12447_));
 sky130_fd_sc_hd__nand3b_4 _35011_ (.A_N(_12446_),
    .B(_12447_),
    .C(_10941_),
    .Y(_12448_));
 sky130_fd_sc_hd__a22o_2 _35012_ (.A1(_10610_),
    .A2(_07004_),
    .B1(_08592_),
    .B2(_07003_),
    .X(_12449_));
 sky130_fd_sc_hd__nand3_2 _35013_ (.A(_12448_),
    .B(_12449_),
    .C(_12442_),
    .Y(_12450_));
 sky130_fd_sc_hd__nand3_4 _35014_ (.A(_12444_),
    .B(_12445_),
    .C(_12450_),
    .Y(_12451_));
 sky130_fd_sc_hd__o21ai_2 _35015_ (.A1(_12440_),
    .A2(_12441_),
    .B1(_12442_),
    .Y(_12452_));
 sky130_fd_sc_hd__nand3_2 _35016_ (.A(_12448_),
    .B(_12449_),
    .C(_12443_),
    .Y(_12453_));
 sky130_fd_sc_hd__o21ai_2 _35017_ (.A1(_12204_),
    .A2(_12202_),
    .B1(_12209_),
    .Y(_12454_));
 sky130_fd_sc_hd__nand3_4 _35018_ (.A(_12452_),
    .B(_12453_),
    .C(_12454_),
    .Y(_12455_));
 sky130_fd_sc_hd__a22oi_4 _35019_ (.A1(_19870_),
    .A2(_07543_),
    .B1(_07902_),
    .B2(_09443_),
    .Y(_12456_));
 sky130_fd_sc_hd__and4_2 _35020_ (.A(_10628_),
    .B(_07973_),
    .C(_07567_),
    .D(_07709_),
    .X(_12457_));
 sky130_fd_sc_hd__nand2_4 _35021_ (.A(_07356_),
    .B(_08042_),
    .Y(_12458_));
 sky130_vsdinv _35022_ (.A(_12458_),
    .Y(_12459_));
 sky130_fd_sc_hd__o21ai_2 _35023_ (.A1(_12456_),
    .A2(_12457_),
    .B1(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__nand2_1 _35024_ (.A(_10628_),
    .B(_07709_),
    .Y(_12461_));
 sky130_fd_sc_hd__nand3b_4 _35025_ (.A_N(_12461_),
    .B(_11871_),
    .C(_10694_),
    .Y(_12462_));
 sky130_fd_sc_hd__a22o_2 _35026_ (.A1(_10934_),
    .A2(_20126_),
    .B1(_10944_),
    .B2(_06976_),
    .X(_12463_));
 sky130_fd_sc_hd__nand3_2 _35027_ (.A(_12462_),
    .B(_12458_),
    .C(_12463_),
    .Y(_12464_));
 sky130_fd_sc_hd__nand2_4 _35028_ (.A(_12460_),
    .B(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__a21o_1 _35029_ (.A1(_12451_),
    .A2(_12455_),
    .B1(_12465_),
    .X(_12466_));
 sky130_fd_sc_hd__nand2_1 _35030_ (.A(_12182_),
    .B(_12187_),
    .Y(_12467_));
 sky130_fd_sc_hd__nand2_2 _35031_ (.A(_12467_),
    .B(_12186_),
    .Y(_12468_));
 sky130_fd_sc_hd__nand3_4 _35032_ (.A(_12451_),
    .B(_12455_),
    .C(_12465_),
    .Y(_12469_));
 sky130_fd_sc_hd__nand3_4 _35033_ (.A(_12466_),
    .B(_12468_),
    .C(_12469_),
    .Y(_12470_));
 sky130_fd_sc_hd__nand2_1 _35034_ (.A(_12466_),
    .B(_12469_),
    .Y(_12471_));
 sky130_fd_sc_hd__a21boi_4 _35035_ (.A1(_12182_),
    .A2(_12187_),
    .B1_N(_12186_),
    .Y(_12472_));
 sky130_fd_sc_hd__and2_1 _35036_ (.A(_12231_),
    .B(_12216_),
    .X(_12473_));
 sky130_fd_sc_hd__a21oi_4 _35037_ (.A1(_12471_),
    .A2(_12472_),
    .B1(_12473_),
    .Y(_12474_));
 sky130_fd_sc_hd__a21oi_4 _35038_ (.A1(_12451_),
    .A2(_12455_),
    .B1(_12465_),
    .Y(_12475_));
 sky130_fd_sc_hd__a21oi_2 _35039_ (.A1(_12462_),
    .A2(_12463_),
    .B1(_12458_),
    .Y(_12476_));
 sky130_fd_sc_hd__and3_1 _35040_ (.A(_12462_),
    .B(_12458_),
    .C(_12463_),
    .X(_12477_));
 sky130_fd_sc_hd__o211a_2 _35041_ (.A1(_12476_),
    .A2(_12477_),
    .B1(_12455_),
    .C1(_12451_),
    .X(_12478_));
 sky130_fd_sc_hd__o21ai_4 _35042_ (.A1(_12475_),
    .A2(_12478_),
    .B1(_12472_),
    .Y(_12479_));
 sky130_fd_sc_hd__nand2_4 _35043_ (.A(_12231_),
    .B(_12216_),
    .Y(_12480_));
 sky130_fd_sc_hd__a21oi_4 _35044_ (.A1(_12479_),
    .A2(_12470_),
    .B1(_12480_),
    .Y(_12481_));
 sky130_fd_sc_hd__a21oi_4 _35045_ (.A1(_12470_),
    .A2(_12474_),
    .B1(_12481_),
    .Y(_12482_));
 sky130_fd_sc_hd__nand2_1 _35046_ (.A(_12146_),
    .B(_12160_),
    .Y(_12483_));
 sky130_fd_sc_hd__nand2_1 _35047_ (.A(_12483_),
    .B(_12150_),
    .Y(_12484_));
 sky130_fd_sc_hd__nand3_4 _35048_ (.A(\pcpi_mul.rs2[32] ),
    .B(\pcpi_mul.rs2[31] ),
    .C(_05480_),
    .Y(_12485_));
 sky130_fd_sc_hd__nor2_8 _35049_ (.A(_06199_),
    .B(_12485_),
    .Y(_12486_));
 sky130_fd_sc_hd__buf_6 _35050_ (.A(_10961_),
    .X(_12487_));
 sky130_fd_sc_hd__a22oi_4 _35051_ (.A1(_10972_),
    .A2(_05481_),
    .B1(_05253_),
    .B2(_12487_),
    .Y(_12488_));
 sky130_fd_sc_hd__nand2_4 _35052_ (.A(_19832_),
    .B(_07417_),
    .Y(_12489_));
 sky130_vsdinv _35053_ (.A(_12489_),
    .Y(_12490_));
 sky130_fd_sc_hd__o21ai_2 _35054_ (.A1(_12486_),
    .A2(_12488_),
    .B1(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__buf_6 _35055_ (.A(_19828_),
    .X(_12492_));
 sky130_fd_sc_hd__o2bb2ai_4 _35056_ (.A1_N(_12492_),
    .A2_N(_06348_),
    .B1(_05238_),
    .B2(_10968_),
    .Y(_12493_));
 sky130_fd_sc_hd__o211ai_4 _35057_ (.A1(_20166_),
    .A2(_12485_),
    .B1(_12489_),
    .C1(_12493_),
    .Y(_12494_));
 sky130_fd_sc_hd__o21ai_1 _35058_ (.A1(_05183_),
    .A2(_12136_),
    .B1(_12139_),
    .Y(_12495_));
 sky130_fd_sc_hd__nand2_2 _35059_ (.A(_12495_),
    .B(_12142_),
    .Y(_12496_));
 sky130_fd_sc_hd__nand3_4 _35060_ (.A(_12491_),
    .B(_12494_),
    .C(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__o21ai_2 _35061_ (.A1(_12486_),
    .A2(_12488_),
    .B1(_12489_),
    .Y(_12498_));
 sky130_fd_sc_hd__nand3b_4 _35062_ (.A_N(_12486_),
    .B(_12490_),
    .C(_12493_),
    .Y(_12499_));
 sky130_fd_sc_hd__o21bai_2 _35063_ (.A1(_12139_),
    .A2(_12138_),
    .B1_N(_12137_),
    .Y(_12500_));
 sky130_fd_sc_hd__nand3_4 _35064_ (.A(_12498_),
    .B(_12499_),
    .C(_12500_),
    .Y(_12501_));
 sky130_fd_sc_hd__nand2_2 _35065_ (.A(_09696_),
    .B(_05699_),
    .Y(_12502_));
 sky130_vsdinv _35066_ (.A(_12502_),
    .Y(_12503_));
 sky130_fd_sc_hd__a22oi_4 _35067_ (.A1(_11794_),
    .A2(_06473_),
    .B1(_19840_),
    .B2(_06476_),
    .Y(_12504_));
 sky130_fd_sc_hd__nand2_2 _35068_ (.A(_09996_),
    .B(_05472_),
    .Y(_12505_));
 sky130_fd_sc_hd__nand2_2 _35069_ (.A(_10989_),
    .B(_05831_),
    .Y(_12506_));
 sky130_fd_sc_hd__nor2_4 _35070_ (.A(_12505_),
    .B(_12506_),
    .Y(_12507_));
 sky130_fd_sc_hd__nor2_1 _35071_ (.A(_12504_),
    .B(_12507_),
    .Y(_12508_));
 sky130_fd_sc_hd__nor2_1 _35072_ (.A(_12503_),
    .B(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__nand3b_4 _35073_ (.A_N(_12505_),
    .B(_09998_),
    .C(_05979_),
    .Y(_12510_));
 sky130_fd_sc_hd__nand2_2 _35074_ (.A(_12505_),
    .B(_12506_),
    .Y(_12511_));
 sky130_fd_sc_hd__and3_1 _35075_ (.A(_12510_),
    .B(_12503_),
    .C(_12511_),
    .X(_12512_));
 sky130_fd_sc_hd__o2bb2ai_2 _35076_ (.A1_N(_12497_),
    .A2_N(_12501_),
    .B1(_12509_),
    .B2(_12512_),
    .Y(_12513_));
 sky130_fd_sc_hd__o21ai_1 _35077_ (.A1(_12504_),
    .A2(_12507_),
    .B1(_12503_),
    .Y(_12514_));
 sky130_fd_sc_hd__nand3_2 _35078_ (.A(_12510_),
    .B(_12502_),
    .C(_12511_),
    .Y(_12515_));
 sky130_fd_sc_hd__nand2_2 _35079_ (.A(_12514_),
    .B(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__nand3_2 _35080_ (.A(_12501_),
    .B(_12497_),
    .C(_12516_),
    .Y(_12517_));
 sky130_fd_sc_hd__nand3_4 _35081_ (.A(_12484_),
    .B(_12513_),
    .C(_12517_),
    .Y(_12518_));
 sky130_vsdinv _35082_ (.A(_12514_),
    .Y(_12519_));
 sky130_vsdinv _35083_ (.A(_12515_),
    .Y(_12520_));
 sky130_fd_sc_hd__o2bb2ai_2 _35084_ (.A1_N(_12497_),
    .A2_N(_12501_),
    .B1(_12519_),
    .B2(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__o21ai_2 _35085_ (.A1(_20169_),
    .A2(_12136_),
    .B1(_12142_),
    .Y(_12522_));
 sky130_fd_sc_hd__a21oi_4 _35086_ (.A1(_12522_),
    .A2(_12139_),
    .B1(_12145_),
    .Y(_12523_));
 sky130_fd_sc_hd__a22oi_4 _35087_ (.A1(_12523_),
    .A2(_12148_),
    .B1(_12146_),
    .B2(_12160_),
    .Y(_12524_));
 sky130_fd_sc_hd__nand3b_2 _35088_ (.A_N(_12516_),
    .B(_12501_),
    .C(_12497_),
    .Y(_12525_));
 sky130_fd_sc_hd__nand3_4 _35089_ (.A(_12521_),
    .B(_12524_),
    .C(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__nand2_2 _35090_ (.A(_12518_),
    .B(_12526_),
    .Y(_12527_));
 sky130_fd_sc_hd__a22oi_4 _35091_ (.A1(_11826_),
    .A2(_20146_),
    .B1(_19851_),
    .B2(_08530_),
    .Y(_12528_));
 sky130_fd_sc_hd__nand3_4 _35092_ (.A(_11008_),
    .B(_09981_),
    .C(_07033_),
    .Y(_12529_));
 sky130_fd_sc_hd__nor2_4 _35093_ (.A(_06307_),
    .B(_12529_),
    .Y(_12530_));
 sky130_fd_sc_hd__nand2_2 _35094_ (.A(_19853_),
    .B(_07502_),
    .Y(_12531_));
 sky130_fd_sc_hd__o21ai_2 _35095_ (.A1(_12528_),
    .A2(_12530_),
    .B1(_12531_),
    .Y(_12532_));
 sky130_vsdinv _35096_ (.A(_12531_),
    .Y(_12533_));
 sky130_fd_sc_hd__a22o_2 _35097_ (.A1(_11826_),
    .A2(_20146_),
    .B1(_19851_),
    .B2(_08530_),
    .X(_12534_));
 sky130_fd_sc_hd__o211ai_4 _35098_ (.A1(_05813_),
    .A2(_12529_),
    .B1(_12533_),
    .C1(_12534_),
    .Y(_12535_));
 sky130_fd_sc_hd__o22ai_4 _35099_ (.A1(net440),
    .A2(_12152_),
    .B1(_12154_),
    .B2(_12157_),
    .Y(_12536_));
 sky130_fd_sc_hd__nand3_4 _35100_ (.A(_12532_),
    .B(_12535_),
    .C(_12536_),
    .Y(_12537_));
 sky130_fd_sc_hd__o21ai_4 _35101_ (.A1(_12528_),
    .A2(_12530_),
    .B1(_12533_),
    .Y(_12538_));
 sky130_fd_sc_hd__a21oi_4 _35102_ (.A1(_12155_),
    .A2(_12158_),
    .B1(_12153_),
    .Y(_12539_));
 sky130_fd_sc_hd__o211ai_4 _35103_ (.A1(_06308_),
    .A2(_12529_),
    .B1(_12531_),
    .C1(_12534_),
    .Y(_12540_));
 sky130_fd_sc_hd__a21oi_4 _35104_ (.A1(_12180_),
    .A2(_12177_),
    .B1(_12175_),
    .Y(_12541_));
 sky130_fd_sc_hd__a31oi_4 _35105_ (.A1(_12538_),
    .A2(_12539_),
    .A3(_12540_),
    .B1(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__nand3_4 _35106_ (.A(_12538_),
    .B(_12539_),
    .C(_12540_),
    .Y(_12543_));
 sky130_vsdinv _35107_ (.A(_12541_),
    .Y(_12544_));
 sky130_fd_sc_hd__a21oi_4 _35108_ (.A1(_12543_),
    .A2(_12537_),
    .B1(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__a21oi_4 _35109_ (.A1(_12537_),
    .A2(_12542_),
    .B1(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__nand2_1 _35110_ (.A(_12527_),
    .B(_12546_),
    .Y(_12547_));
 sky130_fd_sc_hd__a22oi_4 _35111_ (.A1(_11793_),
    .A2(_12169_),
    .B1(_12161_),
    .B2(_12166_),
    .Y(_12548_));
 sky130_fd_sc_hd__a21oi_2 _35112_ (.A1(_12167_),
    .A2(_12193_),
    .B1(_12548_),
    .Y(_12549_));
 sky130_fd_sc_hd__nand3b_2 _35113_ (.A_N(_12546_),
    .B(_12526_),
    .C(_12518_),
    .Y(_12550_));
 sky130_fd_sc_hd__nand3_4 _35114_ (.A(_12547_),
    .B(_12549_),
    .C(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__nand2_2 _35115_ (.A(_12167_),
    .B(_12193_),
    .Y(_12552_));
 sky130_fd_sc_hd__nand2_2 _35116_ (.A(_12552_),
    .B(_12172_),
    .Y(_12553_));
 sky130_fd_sc_hd__and3_1 _35117_ (.A(_12543_),
    .B(_12537_),
    .C(_12544_),
    .X(_12554_));
 sky130_fd_sc_hd__o2bb2ai_2 _35118_ (.A1_N(_12526_),
    .A2_N(_12518_),
    .B1(_12554_),
    .B2(_12545_),
    .Y(_12555_));
 sky130_fd_sc_hd__nand3_4 _35119_ (.A(_12518_),
    .B(_12526_),
    .C(_12546_),
    .Y(_12556_));
 sky130_fd_sc_hd__nand3_4 _35120_ (.A(_12553_),
    .B(_12555_),
    .C(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__nand3_2 _35121_ (.A(_12482_),
    .B(_12551_),
    .C(_12557_),
    .Y(_12558_));
 sky130_fd_sc_hd__nor3_4 _35122_ (.A(_12475_),
    .B(_12472_),
    .C(_12478_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand2_4 _35123_ (.A(_12479_),
    .B(_12480_),
    .Y(_12560_));
 sky130_fd_sc_hd__nor2_1 _35124_ (.A(_12559_),
    .B(_12560_),
    .Y(_12561_));
 sky130_fd_sc_hd__o2bb2ai_2 _35125_ (.A1_N(_12557_),
    .A2_N(_12551_),
    .B1(_12561_),
    .B2(_12481_),
    .Y(_12562_));
 sky130_fd_sc_hd__o211ai_4 _35126_ (.A1(_12254_),
    .A2(_12439_),
    .B1(_12558_),
    .C1(_12562_),
    .Y(_12563_));
 sky130_fd_sc_hd__a21o_1 _35127_ (.A1(_12479_),
    .A2(_12470_),
    .B1(_12480_),
    .X(_12564_));
 sky130_fd_sc_hd__o21ai_4 _35128_ (.A1(_12559_),
    .A2(_12560_),
    .B1(_12564_),
    .Y(_12565_));
 sky130_fd_sc_hd__a21o_1 _35129_ (.A1(_12551_),
    .A2(_12557_),
    .B1(_12565_),
    .X(_12566_));
 sky130_fd_sc_hd__a22oi_4 _35130_ (.A1(_12134_),
    .A2(_11820_),
    .B1(_12196_),
    .B2(_12199_),
    .Y(_12567_));
 sky130_fd_sc_hd__a22oi_4 _35131_ (.A1(_12567_),
    .A2(_12194_),
    .B1(_12201_),
    .B2(_12248_),
    .Y(_12568_));
 sky130_fd_sc_hd__nand3_2 _35132_ (.A(_12565_),
    .B(_12551_),
    .C(_12557_),
    .Y(_12569_));
 sky130_fd_sc_hd__nand3_4 _35133_ (.A(_12566_),
    .B(_12568_),
    .C(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__a22oi_4 _35134_ (.A1(_07088_),
    .A2(_07564_),
    .B1(_07090_),
    .B2(_08056_),
    .Y(_12571_));
 sky130_fd_sc_hd__and4_1 _35135_ (.A(_10067_),
    .B(_06637_),
    .C(_20110_),
    .D(_07233_),
    .X(_12572_));
 sky130_fd_sc_hd__nand2_4 _35136_ (.A(_06640_),
    .B(_08057_),
    .Y(_12573_));
 sky130_fd_sc_hd__o21ai_2 _35137_ (.A1(_12571_),
    .A2(_12572_),
    .B1(_12573_),
    .Y(_12574_));
 sky130_fd_sc_hd__nand2_1 _35138_ (.A(_07294_),
    .B(_08433_),
    .Y(_12575_));
 sky130_fd_sc_hd__buf_6 _35139_ (.A(_07755_),
    .X(_12576_));
 sky130_fd_sc_hd__nand3b_4 _35140_ (.A_N(_12575_),
    .B(_12576_),
    .C(_07723_),
    .Y(_12577_));
 sky130_vsdinv _35141_ (.A(_12573_),
    .Y(_12578_));
 sky130_fd_sc_hd__a22o_1 _35142_ (.A1(_07088_),
    .A2(_07564_),
    .B1(_07449_),
    .B2(_08053_),
    .X(_12579_));
 sky130_fd_sc_hd__nand3_4 _35143_ (.A(_12577_),
    .B(_12578_),
    .C(_12579_),
    .Y(_12580_));
 sky130_fd_sc_hd__o22ai_4 _35144_ (.A1(_08144_),
    .A2(_12219_),
    .B1(_12222_),
    .B2(_12218_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand3_4 _35145_ (.A(_12574_),
    .B(_12580_),
    .C(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__o21ai_2 _35146_ (.A1(_12571_),
    .A2(_12572_),
    .B1(_12578_),
    .Y(_12583_));
 sky130_fd_sc_hd__o22a_1 _35147_ (.A1(_08144_),
    .A2(_12219_),
    .B1(_12222_),
    .B2(_12218_),
    .X(_12584_));
 sky130_fd_sc_hd__nand3_2 _35148_ (.A(_12577_),
    .B(_12573_),
    .C(_12579_),
    .Y(_12585_));
 sky130_fd_sc_hd__nand3_4 _35149_ (.A(_12583_),
    .B(_12584_),
    .C(_12585_),
    .Y(_12586_));
 sky130_fd_sc_hd__nor2_8 _35150_ (.A(_12065_),
    .B(_12062_),
    .Y(_12587_));
 sky130_fd_sc_hd__o2bb2ai_4 _35151_ (.A1_N(_12582_),
    .A2_N(_12586_),
    .B1(_12060_),
    .B2(_12587_),
    .Y(_12588_));
 sky130_fd_sc_hd__nor2_4 _35152_ (.A(_12060_),
    .B(_12587_),
    .Y(_12589_));
 sky130_fd_sc_hd__nand3_4 _35153_ (.A(_12586_),
    .B(_12582_),
    .C(_12589_),
    .Y(_12590_));
 sky130_fd_sc_hd__nand2_1 _35154_ (.A(_12075_),
    .B(_12077_),
    .Y(_12591_));
 sky130_fd_sc_hd__nand2_4 _35155_ (.A(_12591_),
    .B(_12069_),
    .Y(_12592_));
 sky130_fd_sc_hd__a21oi_4 _35156_ (.A1(_12588_),
    .A2(_12590_),
    .B1(_12592_),
    .Y(_12593_));
 sky130_fd_sc_hd__and3_2 _35157_ (.A(_12574_),
    .B(_12580_),
    .C(_12581_),
    .X(_12594_));
 sky130_fd_sc_hd__nand2_2 _35158_ (.A(_12586_),
    .B(_12589_),
    .Y(_12595_));
 sky130_fd_sc_hd__o211a_2 _35159_ (.A1(_12594_),
    .A2(_12595_),
    .B1(_12588_),
    .C1(_12592_),
    .X(_12596_));
 sky130_fd_sc_hd__nor2_4 _35160_ (.A(_12090_),
    .B(_12095_),
    .Y(_12597_));
 sky130_fd_sc_hd__nor2_8 _35161_ (.A(_12088_),
    .B(_12597_),
    .Y(_12598_));
 sky130_fd_sc_hd__a22oi_4 _35162_ (.A1(_06358_),
    .A2(_20105_),
    .B1(_06360_),
    .B2(_09044_),
    .Y(_12599_));
 sky130_fd_sc_hd__nand3_4 _35163_ (.A(_19893_),
    .B(_06359_),
    .C(_20104_),
    .Y(_12600_));
 sky130_fd_sc_hd__nor2_4 _35164_ (.A(_09047_),
    .B(_12600_),
    .Y(_12601_));
 sky130_fd_sc_hd__and2_2 _35165_ (.A(_10700_),
    .B(_09041_),
    .X(_12602_));
 sky130_fd_sc_hd__o21bai_4 _35166_ (.A1(_12599_),
    .A2(_12601_),
    .B1_N(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__buf_4 _35167_ (.A(_09047_),
    .X(_12604_));
 sky130_fd_sc_hd__a22o_1 _35168_ (.A1(_11058_),
    .A2(_08450_),
    .B1(_07422_),
    .B2(_08446_),
    .X(_12605_));
 sky130_fd_sc_hd__o211ai_4 _35169_ (.A1(_12604_),
    .A2(_12600_),
    .B1(_12602_),
    .C1(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__nand2_4 _35170_ (.A(_12603_),
    .B(_12606_),
    .Y(_12607_));
 sky130_fd_sc_hd__nor2_8 _35171_ (.A(_12598_),
    .B(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__nand2_2 _35172_ (.A(_12607_),
    .B(_12598_),
    .Y(_12609_));
 sky130_fd_sc_hd__a22oi_4 _35173_ (.A1(_06042_),
    .A2(_12102_),
    .B1(_07333_),
    .B2(_11210_),
    .Y(_12610_));
 sky130_fd_sc_hd__and4_2 _35174_ (.A(_06042_),
    .B(_07333_),
    .C(_20090_),
    .D(_12102_),
    .X(_12611_));
 sky130_fd_sc_hd__nor2_1 _35175_ (.A(_12610_),
    .B(_12611_),
    .Y(_12612_));
 sky130_fd_sc_hd__nand2_4 _35176_ (.A(_19909_),
    .B(_09474_),
    .Y(_12613_));
 sky130_fd_sc_hd__nand2_1 _35177_ (.A(_12612_),
    .B(_12613_),
    .Y(_12614_));
 sky130_vsdinv _35178_ (.A(_12613_),
    .Y(_12615_));
 sky130_fd_sc_hd__o21ai_1 _35179_ (.A1(_12610_),
    .A2(_12611_),
    .B1(_12615_),
    .Y(_12616_));
 sky130_fd_sc_hd__nand2_2 _35180_ (.A(_12614_),
    .B(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__nand2_1 _35181_ (.A(_12609_),
    .B(_12617_),
    .Y(_12618_));
 sky130_fd_sc_hd__a21o_2 _35182_ (.A1(_12089_),
    .A2(_12091_),
    .B1(_12088_),
    .X(_12619_));
 sky130_fd_sc_hd__a21oi_4 _35183_ (.A1(_12603_),
    .A2(_12606_),
    .B1(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__nand2_1 _35184_ (.A(_12612_),
    .B(_12615_),
    .Y(_12621_));
 sky130_fd_sc_hd__o21ai_1 _35185_ (.A1(_12610_),
    .A2(_12611_),
    .B1(_12613_),
    .Y(_12622_));
 sky130_fd_sc_hd__nand2_2 _35186_ (.A(_12621_),
    .B(_12622_),
    .Y(_12623_));
 sky130_fd_sc_hd__o21ai_2 _35187_ (.A1(_12620_),
    .A2(_12608_),
    .B1(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__o21ai_4 _35188_ (.A1(_12608_),
    .A2(_12618_),
    .B1(_12624_),
    .Y(_12625_));
 sky130_fd_sc_hd__o21ai_2 _35189_ (.A1(_12593_),
    .A2(_12596_),
    .B1(_12625_),
    .Y(_12626_));
 sky130_fd_sc_hd__nand2_2 _35190_ (.A(_12437_),
    .B(_12234_),
    .Y(_12627_));
 sky130_fd_sc_hd__a21o_1 _35191_ (.A1(_12588_),
    .A2(_12590_),
    .B1(_12592_),
    .X(_12628_));
 sky130_fd_sc_hd__nor2_2 _35192_ (.A(_12623_),
    .B(_12620_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand3_4 _35193_ (.A(_12619_),
    .B(_12603_),
    .C(_12606_),
    .Y(_12630_));
 sky130_fd_sc_hd__a21oi_2 _35194_ (.A1(_12609_),
    .A2(_12630_),
    .B1(_12617_),
    .Y(_12631_));
 sky130_fd_sc_hd__a21oi_4 _35195_ (.A1(_12629_),
    .A2(_12630_),
    .B1(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__nand3_4 _35196_ (.A(_12592_),
    .B(_12588_),
    .C(_12590_),
    .Y(_12633_));
 sky130_fd_sc_hd__nand3_4 _35197_ (.A(_12628_),
    .B(_12632_),
    .C(_12633_),
    .Y(_12634_));
 sky130_fd_sc_hd__and3_1 _35198_ (.A(_12626_),
    .B(_12627_),
    .C(_12634_),
    .X(_12635_));
 sky130_fd_sc_hd__o21ai_4 _35199_ (.A1(_12593_),
    .A2(_12596_),
    .B1(_12632_),
    .Y(_12636_));
 sky130_fd_sc_hd__nand3_4 _35200_ (.A(_12628_),
    .B(_12625_),
    .C(_12633_),
    .Y(_12637_));
 sky130_fd_sc_hd__a21boi_4 _35201_ (.A1(_12242_),
    .A2(_12244_),
    .B1_N(_12234_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand3_4 _35202_ (.A(_12636_),
    .B(_12637_),
    .C(_12638_),
    .Y(_12639_));
 sky130_fd_sc_hd__nand2_2 _35203_ (.A(_12278_),
    .B(_12086_),
    .Y(_12640_));
 sky130_fd_sc_hd__nand2_1 _35204_ (.A(_12639_),
    .B(_12640_),
    .Y(_12641_));
 sky130_fd_sc_hd__nor2_2 _35205_ (.A(_12635_),
    .B(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__nand3_4 _35206_ (.A(_12626_),
    .B(_12627_),
    .C(_12634_),
    .Y(_12643_));
 sky130_fd_sc_hd__a21oi_4 _35207_ (.A1(_12643_),
    .A2(_12639_),
    .B1(_12640_),
    .Y(_12644_));
 sky130_fd_sc_hd__o2bb2ai_4 _35208_ (.A1_N(_12563_),
    .A2_N(_12570_),
    .B1(_12642_),
    .B2(_12644_),
    .Y(_12645_));
 sky130_fd_sc_hd__a32oi_4 _35209_ (.A1(_12636_),
    .A2(_12638_),
    .A3(_12637_),
    .B1(_12086_),
    .B2(_12278_),
    .Y(_12646_));
 sky130_fd_sc_hd__a21oi_4 _35210_ (.A1(_12643_),
    .A2(_12646_),
    .B1(_12644_),
    .Y(_12647_));
 sky130_fd_sc_hd__nand3_4 _35211_ (.A(_12647_),
    .B(_12570_),
    .C(_12563_),
    .Y(_12648_));
 sky130_fd_sc_hd__nand3_4 _35212_ (.A(_12434_),
    .B(_12645_),
    .C(_12648_),
    .Y(_12649_));
 sky130_fd_sc_hd__a2bb2oi_4 _35213_ (.A1_N(_12263_),
    .A2_N(_12433_),
    .B1(_12269_),
    .B2(_12265_),
    .Y(_12650_));
 sky130_fd_sc_hd__nand2_1 _35214_ (.A(_12570_),
    .B(_12563_),
    .Y(_12651_));
 sky130_fd_sc_hd__nand2_1 _35215_ (.A(_12651_),
    .B(_12647_),
    .Y(_12652_));
 sky130_fd_sc_hd__nand3b_2 _35216_ (.A_N(_12647_),
    .B(_12570_),
    .C(_12563_),
    .Y(_12653_));
 sky130_fd_sc_hd__nand3_4 _35217_ (.A(_12650_),
    .B(_12652_),
    .C(_12653_),
    .Y(_12654_));
 sky130_fd_sc_hd__nand3b_4 _35218_ (.A_N(_05805_),
    .B(_18686_),
    .C(_19938_),
    .Y(_12655_));
 sky130_fd_sc_hd__nand3_4 _35219_ (.A(_11160_),
    .B(_11603_),
    .C(_19926_),
    .Y(_12656_));
 sky130_fd_sc_hd__inv_2 _35220_ (.A(_19920_),
    .Y(_12657_));
 sky130_fd_sc_hd__o2bb2ai_2 _35221_ (.A1_N(_12655_),
    .A2_N(_12656_),
    .B1(_12657_),
    .B2(_11177_),
    .Y(_12658_));
 sky130_fd_sc_hd__nor2_2 _35222_ (.A(_12657_),
    .B(_11177_),
    .Y(_12659_));
 sky130_fd_sc_hd__nand3_4 _35223_ (.A(_12659_),
    .B(_12655_),
    .C(_12656_),
    .Y(_12660_));
 sky130_fd_sc_hd__a21oi_4 _35224_ (.A1(_11161_),
    .A2(_12338_),
    .B1(_12337_),
    .Y(_12661_));
 sky130_fd_sc_hd__a21o_1 _35225_ (.A1(_12658_),
    .A2(_12660_),
    .B1(_12661_),
    .X(_12662_));
 sky130_fd_sc_hd__nand3_4 _35226_ (.A(_12661_),
    .B(_12658_),
    .C(_12660_),
    .Y(_12663_));
 sky130_fd_sc_hd__a21o_1 _35227_ (.A1(_12662_),
    .A2(_12663_),
    .B1(_12356_),
    .X(_12664_));
 sky130_fd_sc_hd__nand3_4 _35228_ (.A(_12662_),
    .B(_12356_),
    .C(_12663_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand2_1 _35229_ (.A(_12664_),
    .B(_12665_),
    .Y(_12666_));
 sky130_fd_sc_hd__nand2_1 _35230_ (.A(_12346_),
    .B(_12356_),
    .Y(_12667_));
 sky130_fd_sc_hd__nand2_2 _35231_ (.A(_12667_),
    .B(_12342_),
    .Y(_12668_));
 sky130_vsdinv _35232_ (.A(_12668_),
    .Y(_12669_));
 sky130_fd_sc_hd__nand2_1 _35233_ (.A(_12666_),
    .B(_12669_),
    .Y(_12670_));
 sky130_fd_sc_hd__nand3_4 _35234_ (.A(_12664_),
    .B(_12668_),
    .C(_12665_),
    .Y(_12671_));
 sky130_fd_sc_hd__a21oi_4 _35235_ (.A1(_11974_),
    .A2(_19929_),
    .B1(_12330_),
    .Y(_12672_));
 sky130_vsdinv _35236_ (.A(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__buf_2 _35237_ (.A(_12673_),
    .X(_12674_));
 sky130_fd_sc_hd__and3_1 _35238_ (.A(_12670_),
    .B(_12671_),
    .C(_12674_),
    .X(_12675_));
 sky130_fd_sc_hd__a21oi_4 _35239_ (.A1(_12670_),
    .A2(_12671_),
    .B1(_12674_),
    .Y(_12676_));
 sky130_fd_sc_hd__nand2_2 _35240_ (.A(_12319_),
    .B(_12321_),
    .Y(_12677_));
 sky130_fd_sc_hd__a22oi_4 _35241_ (.A1(_06096_),
    .A2(_11157_),
    .B1(_11206_),
    .B2(_10761_),
    .Y(_12678_));
 sky130_fd_sc_hd__nor2_4 _35242_ (.A(_11180_),
    .B(_12291_),
    .Y(_12679_));
 sky130_fd_sc_hd__nand2_2 _35243_ (.A(_05866_),
    .B(_11173_),
    .Y(_12680_));
 sky130_vsdinv _35244_ (.A(_12680_),
    .Y(_12681_));
 sky130_fd_sc_hd__o21ai_2 _35245_ (.A1(_12678_),
    .A2(_12679_),
    .B1(_12681_),
    .Y(_12682_));
 sky130_fd_sc_hd__a21oi_4 _35246_ (.A1(_12107_),
    .A2(_12111_),
    .B1(_12105_),
    .Y(_12683_));
 sky130_fd_sc_hd__a22o_2 _35247_ (.A1(_06096_),
    .A2(_11157_),
    .B1(_06098_),
    .B2(_10761_),
    .X(_12684_));
 sky130_fd_sc_hd__o211ai_4 _35248_ (.A1(_11181_),
    .A2(_12291_),
    .B1(_12680_),
    .C1(_12684_),
    .Y(_12685_));
 sky130_fd_sc_hd__nand3_4 _35249_ (.A(_12682_),
    .B(_12683_),
    .C(_12685_),
    .Y(_12686_));
 sky130_fd_sc_hd__nor2_2 _35250_ (.A(_12106_),
    .B(_12110_),
    .Y(_12687_));
 sky130_fd_sc_hd__buf_6 _35251_ (.A(_11180_),
    .X(_12688_));
 sky130_fd_sc_hd__o211ai_4 _35252_ (.A1(_12688_),
    .A2(_12291_),
    .B1(_12681_),
    .C1(_12684_),
    .Y(_12689_));
 sky130_fd_sc_hd__o21ai_2 _35253_ (.A1(_12678_),
    .A2(_12679_),
    .B1(_12680_),
    .Y(_12690_));
 sky130_fd_sc_hd__o211ai_4 _35254_ (.A1(_12105_),
    .A2(_12687_),
    .B1(_12689_),
    .C1(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__nor2_8 _35255_ (.A(_12294_),
    .B(_12292_),
    .Y(_12692_));
 sky130_fd_sc_hd__o2bb2ai_4 _35256_ (.A1_N(_12686_),
    .A2_N(_12691_),
    .B1(_12290_),
    .B2(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__nor2_8 _35257_ (.A(_12290_),
    .B(_12692_),
    .Y(_12694_));
 sky130_fd_sc_hd__nand3_4 _35258_ (.A(_12691_),
    .B(_12686_),
    .C(_12694_),
    .Y(_12695_));
 sky130_fd_sc_hd__nand2_2 _35259_ (.A(_12124_),
    .B(_12097_),
    .Y(_12696_));
 sky130_fd_sc_hd__a21oi_4 _35260_ (.A1(_12693_),
    .A2(_12695_),
    .B1(_12696_),
    .Y(_12697_));
 sky130_fd_sc_hd__o211a_1 _35261_ (.A1(_12123_),
    .A2(_12113_),
    .B1(_12695_),
    .C1(_12693_),
    .X(_12698_));
 sky130_fd_sc_hd__a21bo_1 _35262_ (.A1(_12301_),
    .A2(_12310_),
    .B1_N(_12309_),
    .X(_12699_));
 sky130_fd_sc_hd__o21bai_4 _35263_ (.A1(_12697_),
    .A2(_12698_),
    .B1_N(_12699_),
    .Y(_12700_));
 sky130_fd_sc_hd__a21oi_1 _35264_ (.A1(_12691_),
    .A2(_12686_),
    .B1(_12694_),
    .Y(_12701_));
 sky130_fd_sc_hd__and3_1 _35265_ (.A(_12691_),
    .B(_12686_),
    .C(_12694_),
    .X(_12702_));
 sky130_fd_sc_hd__o21bai_2 _35266_ (.A1(_12701_),
    .A2(_12702_),
    .B1_N(_12696_),
    .Y(_12703_));
 sky130_fd_sc_hd__nand3_4 _35267_ (.A(_12696_),
    .B(_12693_),
    .C(_12695_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand3_4 _35268_ (.A(_12703_),
    .B(_12704_),
    .C(_12699_),
    .Y(_12705_));
 sky130_fd_sc_hd__a22oi_4 _35269_ (.A1(_12318_),
    .A2(_12677_),
    .B1(_12700_),
    .B2(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__nand2_1 _35270_ (.A(_12703_),
    .B(_12699_),
    .Y(_12707_));
 sky130_fd_sc_hd__o21ai_2 _35271_ (.A1(_12321_),
    .A2(_12313_),
    .B1(_12319_),
    .Y(_12708_));
 sky130_fd_sc_hd__o211a_1 _35272_ (.A1(_12698_),
    .A2(_12707_),
    .B1(_12708_),
    .C1(_12700_),
    .X(_12709_));
 sky130_fd_sc_hd__o22ai_4 _35273_ (.A1(_12675_),
    .A2(_12676_),
    .B1(_12706_),
    .B2(_12709_),
    .Y(_12710_));
 sky130_fd_sc_hd__a21oi_2 _35274_ (.A1(_12666_),
    .A2(_12669_),
    .B1(_12672_),
    .Y(_12711_));
 sky130_fd_sc_hd__a21oi_2 _35275_ (.A1(_12671_),
    .A2(_12711_),
    .B1(_12676_),
    .Y(_12712_));
 sky130_vsdinv _35276_ (.A(_12677_),
    .Y(_12713_));
 sky130_fd_sc_hd__o2bb2ai_2 _35277_ (.A1_N(_12705_),
    .A2_N(_12700_),
    .B1(_12313_),
    .B2(_12713_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand3_4 _35278_ (.A(_12700_),
    .B(_12708_),
    .C(_12705_),
    .Y(_12715_));
 sky130_fd_sc_hd__nand3_4 _35279_ (.A(_12712_),
    .B(_12714_),
    .C(_12715_),
    .Y(_12716_));
 sky130_fd_sc_hd__o21ai_4 _35280_ (.A1(_12276_),
    .A2(_12280_),
    .B1(_12128_),
    .Y(_12717_));
 sky130_fd_sc_hd__a21o_1 _35281_ (.A1(_12710_),
    .A2(_12716_),
    .B1(_12717_),
    .X(_12718_));
 sky130_fd_sc_hd__nand3_4 _35282_ (.A(_12717_),
    .B(_12710_),
    .C(_12716_),
    .Y(_12719_));
 sky130_fd_sc_hd__nand2_4 _35283_ (.A(_12376_),
    .B(_12329_),
    .Y(_12720_));
 sky130_fd_sc_hd__a21oi_2 _35284_ (.A1(_12718_),
    .A2(_12719_),
    .B1(_12720_),
    .Y(_12721_));
 sky130_fd_sc_hd__nand3_4 _35285_ (.A(_12718_),
    .B(_12720_),
    .C(_12719_),
    .Y(_12722_));
 sky130_vsdinv _35286_ (.A(_12722_),
    .Y(_12723_));
 sky130_fd_sc_hd__o2bb2ai_2 _35287_ (.A1_N(_12649_),
    .A2_N(_12654_),
    .B1(_12721_),
    .B2(_12723_),
    .Y(_12724_));
 sky130_fd_sc_hd__o211a_2 _35288_ (.A1(_12279_),
    .A2(_12268_),
    .B1(_12716_),
    .C1(_12710_),
    .X(_12725_));
 sky130_fd_sc_hd__nand2_2 _35289_ (.A(_12718_),
    .B(_12720_),
    .Y(_12726_));
 sky130_fd_sc_hd__a21oi_2 _35290_ (.A1(_12710_),
    .A2(_12716_),
    .B1(_12717_),
    .Y(_12727_));
 sky130_fd_sc_hd__o21bai_4 _35291_ (.A1(_12727_),
    .A2(_12725_),
    .B1_N(_12720_),
    .Y(_12728_));
 sky130_fd_sc_hd__o2111ai_4 _35292_ (.A1(_12725_),
    .A2(_12726_),
    .B1(_12728_),
    .C1(_12649_),
    .D1(_12654_),
    .Y(_12729_));
 sky130_vsdinv _35293_ (.A(_12271_),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_1 _35294_ (.A(_12257_),
    .B(_12272_),
    .Y(_12731_));
 sky130_fd_sc_hd__a21o_1 _35295_ (.A1(_12375_),
    .A2(_12378_),
    .B1(_12379_),
    .X(_12732_));
 sky130_fd_sc_hd__nand2_2 _35296_ (.A(_12732_),
    .B(_12381_),
    .Y(_12733_));
 sky130_fd_sc_hd__a21oi_4 _35297_ (.A1(_12257_),
    .A2(_12271_),
    .B1(_12272_),
    .Y(_12734_));
 sky130_fd_sc_hd__o22ai_4 _35298_ (.A1(_12730_),
    .A2(_12731_),
    .B1(_12733_),
    .B2(_12734_),
    .Y(_12735_));
 sky130_fd_sc_hd__a21oi_4 _35299_ (.A1(_12724_),
    .A2(_12729_),
    .B1(_12735_),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_2 _35300_ (.A(_12386_),
    .B(_12284_),
    .Y(_12737_));
 sky130_fd_sc_hd__a22oi_4 _35301_ (.A1(_12728_),
    .A2(_12722_),
    .B1(_12654_),
    .B2(_12649_),
    .Y(_12738_));
 sky130_fd_sc_hd__o2111a_4 _35302_ (.A1(_12725_),
    .A2(_12726_),
    .B1(_12728_),
    .C1(_12649_),
    .D1(_12654_),
    .X(_12739_));
 sky130_fd_sc_hd__a211oi_4 _35303_ (.A1(_12737_),
    .A2(_12273_),
    .B1(_12738_),
    .C1(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__o22ai_4 _35304_ (.A1(_12430_),
    .A2(_12432_),
    .B1(_12736_),
    .B2(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__a21oi_4 _35305_ (.A1(_12737_),
    .A2(_12273_),
    .B1(_12738_),
    .Y(_12742_));
 sky130_fd_sc_hd__nand2_2 _35306_ (.A(_12742_),
    .B(_12729_),
    .Y(_12743_));
 sky130_fd_sc_hd__o21a_1 _35307_ (.A1(_12733_),
    .A2(_12734_),
    .B1(_12273_),
    .X(_12744_));
 sky130_fd_sc_hd__o21ai_4 _35308_ (.A1(_12738_),
    .A2(_12739_),
    .B1(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__nor2_4 _35309_ (.A(_12432_),
    .B(_12430_),
    .Y(_12746_));
 sky130_fd_sc_hd__nand3_4 _35310_ (.A(_12743_),
    .B(_12745_),
    .C(_12746_),
    .Y(_12747_));
 sky130_fd_sc_hd__nand3_4 _35311_ (.A(_12425_),
    .B(_12741_),
    .C(_12747_),
    .Y(_12748_));
 sky130_fd_sc_hd__nor2_8 _35312_ (.A(_12431_),
    .B(_12429_),
    .Y(_12749_));
 sky130_fd_sc_hd__nor2_4 _35313_ (.A(_12427_),
    .B(_12428_),
    .Y(_12750_));
 sky130_fd_sc_hd__o22ai_4 _35314_ (.A1(_12749_),
    .A2(_12750_),
    .B1(_12736_),
    .B2(_12740_),
    .Y(_12751_));
 sky130_fd_sc_hd__nor2_4 _35315_ (.A(_12750_),
    .B(_12749_),
    .Y(_12752_));
 sky130_fd_sc_hd__nand3_4 _35316_ (.A(_12743_),
    .B(_12745_),
    .C(_12752_),
    .Y(_12753_));
 sky130_fd_sc_hd__o21ai_2 _35317_ (.A1(_12401_),
    .A2(_12389_),
    .B1(_12402_),
    .Y(_12754_));
 sky130_fd_sc_hd__nand3_4 _35318_ (.A(_12751_),
    .B(_12753_),
    .C(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__a21oi_4 _35319_ (.A1(_12748_),
    .A2(_12755_),
    .B1(_12405_),
    .Y(_12756_));
 sky130_fd_sc_hd__and3_1 _35320_ (.A(_12748_),
    .B(_12755_),
    .C(_12405_),
    .X(_12757_));
 sky130_vsdinv _35321_ (.A(_12406_),
    .Y(_12758_));
 sky130_fd_sc_hd__nand2_1 _35322_ (.A(_12408_),
    .B(_12407_),
    .Y(_12759_));
 sky130_fd_sc_hd__o2bb2ai_4 _35323_ (.A1_N(_12037_),
    .A2_N(_12404_),
    .B1(_12758_),
    .B2(_12759_),
    .Y(_12760_));
 sky130_fd_sc_hd__o21bai_2 _35324_ (.A1(_12756_),
    .A2(_12757_),
    .B1_N(_12760_),
    .Y(_12761_));
 sky130_fd_sc_hd__a21o_1 _35325_ (.A1(_12748_),
    .A2(_12755_),
    .B1(_12405_),
    .X(_12762_));
 sky130_fd_sc_hd__nand3_4 _35326_ (.A(_12748_),
    .B(_12755_),
    .C(_12405_),
    .Y(_12763_));
 sky130_fd_sc_hd__nand3_4 _35327_ (.A(_12762_),
    .B(_12760_),
    .C(_12763_),
    .Y(_12764_));
 sky130_fd_sc_hd__nand2_1 _35328_ (.A(_12761_),
    .B(_12764_),
    .Y(_12765_));
 sky130_fd_sc_hd__and3_1 _35329_ (.A(_12053_),
    .B(_12052_),
    .C(_12422_),
    .X(_12766_));
 sky130_fd_sc_hd__o2111ai_4 _35330_ (.A1(_12411_),
    .A2(_12417_),
    .B1(_12051_),
    .C1(_12048_),
    .D1(_12421_),
    .Y(_12767_));
 sky130_fd_sc_hd__a21oi_1 _35331_ (.A1(_12418_),
    .A2(_12410_),
    .B1(_12420_),
    .Y(_12768_));
 sky130_fd_sc_hd__o22ai_1 _35332_ (.A1(_12411_),
    .A2(_12417_),
    .B1(_12051_),
    .B2(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__o21bai_4 _35333_ (.A1(_12055_),
    .A2(_12767_),
    .B1_N(_12769_),
    .Y(_12770_));
 sky130_fd_sc_hd__a21oi_4 _35334_ (.A1(net409),
    .A2(_12766_),
    .B1(_12770_),
    .Y(_12771_));
 sky130_fd_sc_hd__or2_1 _35335_ (.A(_12765_),
    .B(_12771_),
    .X(_12772_));
 sky130_fd_sc_hd__nand2_1 _35336_ (.A(_12771_),
    .B(_12765_),
    .Y(_12773_));
 sky130_fd_sc_hd__and2_4 _35337_ (.A(_12772_),
    .B(_12773_),
    .X(_02655_));
 sky130_fd_sc_hd__a21oi_2 _35338_ (.A1(_12555_),
    .A2(_12556_),
    .B1(_12553_),
    .Y(_12774_));
 sky130_fd_sc_hd__o21ai_4 _35339_ (.A1(_12565_),
    .A2(_12774_),
    .B1(_12557_),
    .Y(_12775_));
 sky130_fd_sc_hd__nand3_4 _35340_ (.A(_18693_),
    .B(_19828_),
    .C(_05391_),
    .Y(_12776_));
 sky130_fd_sc_hd__nor2_8 _35341_ (.A(_05867_),
    .B(_12776_),
    .Y(_12777_));
 sky130_fd_sc_hd__a22oi_4 _35342_ (.A1(_12492_),
    .A2(_05675_),
    .B1(_09275_),
    .B2(_12487_),
    .Y(_12778_));
 sky130_fd_sc_hd__nand2_2 _35343_ (.A(_10577_),
    .B(_05981_),
    .Y(_12779_));
 sky130_vsdinv _35344_ (.A(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__o21ai_2 _35345_ (.A1(_12777_),
    .A2(_12778_),
    .B1(_12780_),
    .Y(_12781_));
 sky130_fd_sc_hd__o2bb2ai_4 _35346_ (.A1_N(_12492_),
    .A2_N(_20159_),
    .B1(_06348_),
    .B2(_10968_),
    .Y(_12782_));
 sky130_fd_sc_hd__nand3b_2 _35347_ (.A_N(_12777_),
    .B(_12779_),
    .C(_12782_),
    .Y(_12783_));
 sky130_fd_sc_hd__a21oi_4 _35348_ (.A1(_12493_),
    .A2(_12490_),
    .B1(_12486_),
    .Y(_12784_));
 sky130_fd_sc_hd__nand3_4 _35349_ (.A(_12781_),
    .B(_12783_),
    .C(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__o21ai_2 _35350_ (.A1(_12777_),
    .A2(_12778_),
    .B1(_12779_),
    .Y(_12786_));
 sky130_fd_sc_hd__o211ai_4 _35351_ (.A1(_20163_),
    .A2(_12776_),
    .B1(_12780_),
    .C1(_12782_),
    .Y(_12787_));
 sky130_fd_sc_hd__o22ai_4 _35352_ (.A1(_20166_),
    .A2(_12485_),
    .B1(_12489_),
    .B2(_12488_),
    .Y(_12788_));
 sky130_fd_sc_hd__nand3_4 _35353_ (.A(_12786_),
    .B(_12787_),
    .C(_12788_),
    .Y(_12789_));
 sky130_fd_sc_hd__nor2_8 _35354_ (.A(_05690_),
    .B(_10983_),
    .Y(_12790_));
 sky130_fd_sc_hd__nand2_2 _35355_ (.A(_19843_),
    .B(_05835_),
    .Y(_12791_));
 sky130_fd_sc_hd__a22o_2 _35356_ (.A1(_10411_),
    .A2(_06476_),
    .B1(_10412_),
    .B2(_10611_),
    .X(_12792_));
 sky130_fd_sc_hd__nand3b_4 _35357_ (.A_N(_12790_),
    .B(_12791_),
    .C(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__a22oi_4 _35358_ (.A1(_09997_),
    .A2(_05991_),
    .B1(_09998_),
    .B2(_05820_),
    .Y(_12794_));
 sky130_vsdinv _35359_ (.A(_12791_),
    .Y(_12795_));
 sky130_fd_sc_hd__o21ai_2 _35360_ (.A1(_12794_),
    .A2(_12790_),
    .B1(_12795_),
    .Y(_12796_));
 sky130_fd_sc_hd__nand2_4 _35361_ (.A(_12793_),
    .B(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__a21o_1 _35362_ (.A1(_12785_),
    .A2(_12789_),
    .B1(_12797_),
    .X(_12798_));
 sky130_fd_sc_hd__nand2_1 _35363_ (.A(_12497_),
    .B(_12516_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand2_2 _35364_ (.A(_12799_),
    .B(_12501_),
    .Y(_12800_));
 sky130_fd_sc_hd__nand3_2 _35365_ (.A(_12785_),
    .B(_12789_),
    .C(_12797_),
    .Y(_12801_));
 sky130_fd_sc_hd__nand3_4 _35366_ (.A(_12798_),
    .B(_12800_),
    .C(_12801_),
    .Y(_12802_));
 sky130_vsdinv _35367_ (.A(_12796_),
    .Y(_12803_));
 sky130_vsdinv _35368_ (.A(_12793_),
    .Y(_12804_));
 sky130_fd_sc_hd__o2bb2ai_4 _35369_ (.A1_N(_12789_),
    .A2_N(_12785_),
    .B1(_12803_),
    .B2(_12804_),
    .Y(_12805_));
 sky130_fd_sc_hd__o21ai_1 _35370_ (.A1(_20166_),
    .A2(_12485_),
    .B1(_12493_),
    .Y(_12806_));
 sky130_fd_sc_hd__a21oi_2 _35371_ (.A1(_12806_),
    .A2(_12489_),
    .B1(_12496_),
    .Y(_12807_));
 sky130_fd_sc_hd__a22oi_4 _35372_ (.A1(_12807_),
    .A2(_12499_),
    .B1(_12497_),
    .B2(_12516_),
    .Y(_12808_));
 sky130_fd_sc_hd__nand3b_4 _35373_ (.A_N(_12797_),
    .B(_12785_),
    .C(_12789_),
    .Y(_12809_));
 sky130_fd_sc_hd__nand3_4 _35374_ (.A(_12805_),
    .B(_12808_),
    .C(_12809_),
    .Y(_12810_));
 sky130_fd_sc_hd__a22oi_4 _35375_ (.A1(_11826_),
    .A2(_08530_),
    .B1(_19851_),
    .B2(_06151_),
    .Y(_12811_));
 sky130_fd_sc_hd__nand3_4 _35376_ (.A(_10383_),
    .B(_08800_),
    .C(_06154_),
    .Y(_12812_));
 sky130_fd_sc_hd__nor2_4 _35377_ (.A(net465),
    .B(_12812_),
    .Y(_12813_));
 sky130_fd_sc_hd__nand2_4 _35378_ (.A(_19854_),
    .B(_06312_),
    .Y(_12814_));
 sky130_vsdinv _35379_ (.A(_12814_),
    .Y(_12815_));
 sky130_fd_sc_hd__o21ai_2 _35380_ (.A1(_12811_),
    .A2(_12813_),
    .B1(_12815_),
    .Y(_12816_));
 sky130_fd_sc_hd__a21oi_4 _35381_ (.A1(_12503_),
    .A2(_12511_),
    .B1(_12507_),
    .Y(_12817_));
 sky130_fd_sc_hd__buf_4 _35382_ (.A(_08800_),
    .X(_12818_));
 sky130_fd_sc_hd__a22o_2 _35383_ (.A1(_11366_),
    .A2(_20143_),
    .B1(_12818_),
    .B2(net466),
    .X(_12819_));
 sky130_fd_sc_hd__o211ai_4 _35384_ (.A1(_07191_),
    .A2(_12812_),
    .B1(_12814_),
    .C1(_12819_),
    .Y(_12820_));
 sky130_fd_sc_hd__nand3_4 _35385_ (.A(_12816_),
    .B(_12817_),
    .C(_12820_),
    .Y(_12821_));
 sky130_fd_sc_hd__o21ai_2 _35386_ (.A1(_12811_),
    .A2(_12813_),
    .B1(_12814_),
    .Y(_12822_));
 sky130_fd_sc_hd__o21ai_2 _35387_ (.A1(_12502_),
    .A2(_12504_),
    .B1(_12510_),
    .Y(_12823_));
 sky130_fd_sc_hd__o211ai_4 _35388_ (.A1(_07191_),
    .A2(_12812_),
    .B1(_12815_),
    .C1(_12819_),
    .Y(_12824_));
 sky130_fd_sc_hd__nand3_4 _35389_ (.A(_12822_),
    .B(_12823_),
    .C(_12824_),
    .Y(_12825_));
 sky130_fd_sc_hd__nor2_2 _35390_ (.A(_12533_),
    .B(_12530_),
    .Y(_12826_));
 sky130_fd_sc_hd__o2bb2ai_2 _35391_ (.A1_N(_12821_),
    .A2_N(_12825_),
    .B1(_12528_),
    .B2(_12826_),
    .Y(_12827_));
 sky130_fd_sc_hd__nor2_2 _35392_ (.A(_12528_),
    .B(_12826_),
    .Y(_12828_));
 sky130_fd_sc_hd__nand3_2 _35393_ (.A(_12821_),
    .B(_12825_),
    .C(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__nand2_2 _35394_ (.A(_12827_),
    .B(_12829_),
    .Y(_12830_));
 sky130_fd_sc_hd__a21o_1 _35395_ (.A1(_12802_),
    .A2(_12810_),
    .B1(_12830_),
    .X(_12831_));
 sky130_fd_sc_hd__a21boi_2 _35396_ (.A1(_12526_),
    .A2(_12546_),
    .B1_N(_12518_),
    .Y(_12832_));
 sky130_fd_sc_hd__nand3_2 _35397_ (.A(_12802_),
    .B(_12810_),
    .C(_12830_),
    .Y(_12833_));
 sky130_fd_sc_hd__nand3_4 _35398_ (.A(_12831_),
    .B(_12832_),
    .C(_12833_),
    .Y(_12834_));
 sky130_fd_sc_hd__nand2_1 _35399_ (.A(_12526_),
    .B(_12546_),
    .Y(_12835_));
 sky130_fd_sc_hd__nand2_2 _35400_ (.A(_12835_),
    .B(_12518_),
    .Y(_12836_));
 sky130_vsdinv _35401_ (.A(_12827_),
    .Y(_12837_));
 sky130_vsdinv _35402_ (.A(_12829_),
    .Y(_12838_));
 sky130_fd_sc_hd__o2bb2ai_2 _35403_ (.A1_N(_12810_),
    .A2_N(_12802_),
    .B1(_12837_),
    .B2(_12838_),
    .Y(_12839_));
 sky130_vsdinv _35404_ (.A(_12825_),
    .Y(_12840_));
 sky130_fd_sc_hd__nand2_2 _35405_ (.A(_12821_),
    .B(_12828_),
    .Y(_12841_));
 sky130_fd_sc_hd__o21a_2 _35406_ (.A1(_12840_),
    .A2(_12841_),
    .B1(_12827_),
    .X(_12842_));
 sky130_fd_sc_hd__nand3_4 _35407_ (.A(_12802_),
    .B(_12842_),
    .C(_12810_),
    .Y(_12843_));
 sky130_fd_sc_hd__nand3_4 _35408_ (.A(_12836_),
    .B(_12839_),
    .C(_12843_),
    .Y(_12844_));
 sky130_fd_sc_hd__nand2_2 _35409_ (.A(_12537_),
    .B(_12541_),
    .Y(_12845_));
 sky130_fd_sc_hd__buf_6 _35410_ (.A(_08151_),
    .X(_12846_));
 sky130_fd_sc_hd__a22oi_4 _35411_ (.A1(_19859_),
    .A2(_20134_),
    .B1(_10918_),
    .B2(_12846_),
    .Y(_12847_));
 sky130_fd_sc_hd__clkbuf_4 _35412_ (.A(_19858_),
    .X(_12848_));
 sky130_fd_sc_hd__and4_2 _35413_ (.A(_12848_),
    .B(_19863_),
    .C(_20130_),
    .D(_08546_),
    .X(_12849_));
 sky130_fd_sc_hd__nand2_2 _35414_ (.A(_07967_),
    .B(_07543_),
    .Y(_12850_));
 sky130_vsdinv _35415_ (.A(_12850_),
    .Y(_12851_));
 sky130_fd_sc_hd__o21ai_2 _35416_ (.A1(_12847_),
    .A2(_12849_),
    .B1(_12851_),
    .Y(_12852_));
 sky130_fd_sc_hd__a21oi_4 _35417_ (.A1(_12449_),
    .A2(_12443_),
    .B1(_12441_),
    .Y(_12853_));
 sky130_fd_sc_hd__nand2_1 _35418_ (.A(_12848_),
    .B(_08546_),
    .Y(_12854_));
 sky130_fd_sc_hd__buf_4 _35419_ (.A(_08592_),
    .X(_12855_));
 sky130_fd_sc_hd__nand3b_4 _35420_ (.A_N(_12854_),
    .B(_12855_),
    .C(_12846_),
    .Y(_12856_));
 sky130_fd_sc_hd__a22o_2 _35421_ (.A1(_10917_),
    .A2(_10941_),
    .B1(_12447_),
    .B2(_11093_),
    .X(_12857_));
 sky130_fd_sc_hd__nand3_2 _35422_ (.A(_12856_),
    .B(_12857_),
    .C(_12850_),
    .Y(_12858_));
 sky130_fd_sc_hd__nand3_4 _35423_ (.A(_12852_),
    .B(_12853_),
    .C(_12858_),
    .Y(_12859_));
 sky130_fd_sc_hd__o21ai_2 _35424_ (.A1(_12847_),
    .A2(_12849_),
    .B1(_12850_),
    .Y(_12860_));
 sky130_fd_sc_hd__nand3_2 _35425_ (.A(_12856_),
    .B(_12857_),
    .C(_12851_),
    .Y(_12861_));
 sky130_fd_sc_hd__o21ai_2 _35426_ (.A1(_12442_),
    .A2(_12440_),
    .B1(_12448_),
    .Y(_12862_));
 sky130_fd_sc_hd__nand3_4 _35427_ (.A(_12860_),
    .B(_12861_),
    .C(_12862_),
    .Y(_12863_));
 sky130_fd_sc_hd__buf_4 _35428_ (.A(_08326_),
    .X(_12864_));
 sky130_fd_sc_hd__a22oi_4 _35429_ (.A1(_12864_),
    .A2(_09443_),
    .B1(_11871_),
    .B2(_12059_),
    .Y(_12865_));
 sky130_fd_sc_hd__and4_2 _35430_ (.A(_12864_),
    .B(_11871_),
    .C(_07726_),
    .D(_10694_),
    .X(_12866_));
 sky130_fd_sc_hd__nor2_1 _35431_ (.A(_12865_),
    .B(_12866_),
    .Y(_12867_));
 sky130_fd_sc_hd__nand2_2 _35432_ (.A(_11869_),
    .B(_08060_),
    .Y(_12868_));
 sky130_fd_sc_hd__nand2_1 _35433_ (.A(_12867_),
    .B(_12868_),
    .Y(_12869_));
 sky130_vsdinv _35434_ (.A(_12868_),
    .Y(_12870_));
 sky130_fd_sc_hd__o21ai_1 _35435_ (.A1(_12865_),
    .A2(_12866_),
    .B1(_12870_),
    .Y(_12871_));
 sky130_fd_sc_hd__nand2_2 _35436_ (.A(_12869_),
    .B(_12871_),
    .Y(_12872_));
 sky130_fd_sc_hd__a21oi_2 _35437_ (.A1(_12859_),
    .A2(_12863_),
    .B1(_12872_),
    .Y(_12873_));
 sky130_fd_sc_hd__nor3_2 _35438_ (.A(_12870_),
    .B(_12865_),
    .C(_12866_),
    .Y(_12874_));
 sky130_fd_sc_hd__o21a_1 _35439_ (.A1(_12865_),
    .A2(_12866_),
    .B1(_12870_),
    .X(_12875_));
 sky130_fd_sc_hd__o211a_2 _35440_ (.A1(_12874_),
    .A2(_12875_),
    .B1(_12863_),
    .C1(_12859_),
    .X(_12876_));
 sky130_fd_sc_hd__o2bb2ai_4 _35441_ (.A1_N(_12543_),
    .A2_N(_12845_),
    .B1(_12873_),
    .B2(_12876_),
    .Y(_12877_));
 sky130_fd_sc_hd__and3_1 _35442_ (.A(_12532_),
    .B(_12535_),
    .C(_12536_),
    .X(_12878_));
 sky130_vsdinv _35443_ (.A(_12863_),
    .Y(_12879_));
 sky130_fd_sc_hd__nand2_2 _35444_ (.A(_12872_),
    .B(_12859_),
    .Y(_12880_));
 sky130_fd_sc_hd__a21o_1 _35445_ (.A1(_12859_),
    .A2(_12863_),
    .B1(_12872_),
    .X(_12881_));
 sky130_fd_sc_hd__o221ai_4 _35446_ (.A1(_12878_),
    .A2(_12542_),
    .B1(_12879_),
    .B2(_12880_),
    .C1(_12881_),
    .Y(_12882_));
 sky130_vsdinv _35447_ (.A(_12455_),
    .Y(_12883_));
 sky130_fd_sc_hd__a21o_2 _35448_ (.A1(_12451_),
    .A2(_12465_),
    .B1(_12883_),
    .X(_12884_));
 sky130_fd_sc_hd__a21oi_4 _35449_ (.A1(_12877_),
    .A2(_12882_),
    .B1(_12884_),
    .Y(_12885_));
 sky130_fd_sc_hd__and2_1 _35450_ (.A(_12451_),
    .B(_12465_),
    .X(_12886_));
 sky130_fd_sc_hd__o211a_2 _35451_ (.A1(_12883_),
    .A2(_12886_),
    .B1(_12882_),
    .C1(_12877_),
    .X(_12887_));
 sky130_fd_sc_hd__o2bb2ai_4 _35452_ (.A1_N(_12834_),
    .A2_N(_12844_),
    .B1(_12885_),
    .B2(_12887_),
    .Y(_12888_));
 sky130_fd_sc_hd__nor2_4 _35453_ (.A(_12885_),
    .B(_12887_),
    .Y(_12889_));
 sky130_fd_sc_hd__nand3_4 _35454_ (.A(_12889_),
    .B(_12834_),
    .C(_12844_),
    .Y(_12890_));
 sky130_fd_sc_hd__nand3_4 _35455_ (.A(_12775_),
    .B(_12888_),
    .C(_12890_),
    .Y(_12891_));
 sky130_fd_sc_hd__nand2_1 _35456_ (.A(_12834_),
    .B(_12844_),
    .Y(_12892_));
 sky130_fd_sc_hd__nand2_1 _35457_ (.A(_12892_),
    .B(_12889_),
    .Y(_12893_));
 sky130_vsdinv _35458_ (.A(_12546_),
    .Y(_12894_));
 sky130_fd_sc_hd__a22oi_4 _35459_ (.A1(_12552_),
    .A2(_12172_),
    .B1(_12527_),
    .B2(_12894_),
    .Y(_12895_));
 sky130_fd_sc_hd__a22oi_4 _35460_ (.A1(_12895_),
    .A2(_12556_),
    .B1(_12482_),
    .B2(_12551_),
    .Y(_12896_));
 sky130_fd_sc_hd__a21o_1 _35461_ (.A1(_12877_),
    .A2(_12882_),
    .B1(_12884_),
    .X(_12897_));
 sky130_fd_sc_hd__nand3_2 _35462_ (.A(_12877_),
    .B(_12882_),
    .C(_12884_),
    .Y(_12898_));
 sky130_fd_sc_hd__nand2_1 _35463_ (.A(_12897_),
    .B(_12898_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand3_2 _35464_ (.A(_12899_),
    .B(_12834_),
    .C(_12844_),
    .Y(_12900_));
 sky130_fd_sc_hd__nand3_4 _35465_ (.A(_12893_),
    .B(_12896_),
    .C(_12900_),
    .Y(_12901_));
 sky130_fd_sc_hd__nand2_1 _35466_ (.A(_12891_),
    .B(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__and4_2 _35467_ (.A(_11058_),
    .B(_07422_),
    .C(_09041_),
    .D(_08446_),
    .X(_12903_));
 sky130_fd_sc_hd__a22o_1 _35468_ (.A1(_11486_),
    .A2(_08446_),
    .B1(_07115_),
    .B2(_12103_),
    .X(_12904_));
 sky130_fd_sc_hd__nand2_2 _35469_ (.A(_10700_),
    .B(_20093_),
    .Y(_12905_));
 sky130_vsdinv _35470_ (.A(_12905_),
    .Y(_12906_));
 sky130_fd_sc_hd__nand2_4 _35471_ (.A(_12904_),
    .B(_12906_),
    .Y(_12907_));
 sky130_fd_sc_hd__a22oi_4 _35472_ (.A1(_10692_),
    .A2(_10222_),
    .B1(_10693_),
    .B2(_11503_),
    .Y(_12908_));
 sky130_fd_sc_hd__o21ai_2 _35473_ (.A1(_12908_),
    .A2(_12903_),
    .B1(_12905_),
    .Y(_12909_));
 sky130_fd_sc_hd__a21o_1 _35474_ (.A1(_12605_),
    .A2(_12602_),
    .B1(_12601_),
    .X(_12910_));
 sky130_fd_sc_hd__o211ai_4 _35475_ (.A1(_12903_),
    .A2(_12907_),
    .B1(_12909_),
    .C1(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__o21ai_2 _35476_ (.A1(_12908_),
    .A2(_12903_),
    .B1(_12906_),
    .Y(_12912_));
 sky130_fd_sc_hd__a21oi_2 _35477_ (.A1(_12605_),
    .A2(_12602_),
    .B1(_12601_),
    .Y(_12913_));
 sky130_fd_sc_hd__nand2_1 _35478_ (.A(_11058_),
    .B(_08446_),
    .Y(_12914_));
 sky130_fd_sc_hd__nand3b_4 _35479_ (.A_N(_12914_),
    .B(_06360_),
    .C(_09493_),
    .Y(_12915_));
 sky130_fd_sc_hd__nand3_2 _35480_ (.A(_12915_),
    .B(_12904_),
    .C(_12905_),
    .Y(_12916_));
 sky130_fd_sc_hd__nand3_4 _35481_ (.A(_12912_),
    .B(_12913_),
    .C(_12916_),
    .Y(_12917_));
 sky130_fd_sc_hd__nand2_1 _35482_ (.A(_12911_),
    .B(_12917_),
    .Y(_12918_));
 sky130_fd_sc_hd__a22oi_4 _35483_ (.A1(_19902_),
    .A2(_09487_),
    .B1(_06049_),
    .B2(_09787_),
    .Y(_12919_));
 sky130_fd_sc_hd__nand2_2 _35484_ (.A(_06630_),
    .B(\pcpi_mul.rs1[26] ),
    .Y(_12920_));
 sky130_fd_sc_hd__nand2_2 _35485_ (.A(_06045_),
    .B(_09474_),
    .Y(_12921_));
 sky130_fd_sc_hd__nor2_1 _35486_ (.A(_12920_),
    .B(_12921_),
    .Y(_12922_));
 sky130_fd_sc_hd__nand2_2 _35487_ (.A(_06052_),
    .B(_10259_),
    .Y(_12923_));
 sky130_fd_sc_hd__o21bai_2 _35488_ (.A1(_12919_),
    .A2(_12922_),
    .B1_N(_12923_),
    .Y(_12924_));
 sky130_fd_sc_hd__nand3b_4 _35489_ (.A_N(_12920_),
    .B(_10347_),
    .C(_11934_),
    .Y(_12925_));
 sky130_fd_sc_hd__nand2_1 _35490_ (.A(_12920_),
    .B(_12921_),
    .Y(_12926_));
 sky130_fd_sc_hd__nand3_2 _35491_ (.A(_12925_),
    .B(_12923_),
    .C(_12926_),
    .Y(_12927_));
 sky130_fd_sc_hd__nand2_4 _35492_ (.A(_12924_),
    .B(_12927_),
    .Y(_12928_));
 sky130_fd_sc_hd__and2_1 _35493_ (.A(_12918_),
    .B(_12928_),
    .X(_12929_));
 sky130_fd_sc_hd__nor2_2 _35494_ (.A(_12928_),
    .B(_12918_),
    .Y(_12930_));
 sky130_fd_sc_hd__a22oi_4 _35495_ (.A1(_11092_),
    .A2(_07723_),
    .B1(_19887_),
    .B2(_08453_),
    .Y(_12931_));
 sky130_fd_sc_hd__nand3_4 _35496_ (.A(_10067_),
    .B(_06637_),
    .C(_20110_),
    .Y(_12932_));
 sky130_fd_sc_hd__nor2_4 _35497_ (.A(_09732_),
    .B(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__nand2_2 _35498_ (.A(_19890_),
    .B(_20104_),
    .Y(_12934_));
 sky130_vsdinv _35499_ (.A(_12934_),
    .Y(_12935_));
 sky130_fd_sc_hd__o21ai_2 _35500_ (.A1(_12931_),
    .A2(_12933_),
    .B1(_12935_),
    .Y(_12936_));
 sky130_fd_sc_hd__a21oi_4 _35501_ (.A1(_12463_),
    .A2(_12459_),
    .B1(_12457_),
    .Y(_12937_));
 sky130_fd_sc_hd__a22o_4 _35502_ (.A1(_19881_),
    .A2(_08056_),
    .B1(_12576_),
    .B2(_08052_),
    .X(_12938_));
 sky130_fd_sc_hd__o211ai_4 _35503_ (.A1(_11734_),
    .A2(_12932_),
    .B1(_12934_),
    .C1(_12938_),
    .Y(_12939_));
 sky130_fd_sc_hd__nand3_4 _35504_ (.A(_12936_),
    .B(_12937_),
    .C(_12939_),
    .Y(_12940_));
 sky130_fd_sc_hd__o21ai_2 _35505_ (.A1(_12931_),
    .A2(_12933_),
    .B1(_12934_),
    .Y(_12941_));
 sky130_fd_sc_hd__o211ai_4 _35506_ (.A1(_11734_),
    .A2(_12932_),
    .B1(_12935_),
    .C1(_12938_),
    .Y(_12942_));
 sky130_fd_sc_hd__o21ai_2 _35507_ (.A1(_12458_),
    .A2(_12456_),
    .B1(_12462_),
    .Y(_12943_));
 sky130_fd_sc_hd__nand3_4 _35508_ (.A(_12941_),
    .B(_12942_),
    .C(_12943_),
    .Y(_12944_));
 sky130_fd_sc_hd__o21ai_4 _35509_ (.A1(_12573_),
    .A2(_12571_),
    .B1(_12577_),
    .Y(_12945_));
 sky130_fd_sc_hd__a21o_2 _35510_ (.A1(_12940_),
    .A2(_12944_),
    .B1(_12945_),
    .X(_12946_));
 sky130_fd_sc_hd__nand3_4 _35511_ (.A(_12940_),
    .B(_12944_),
    .C(_12945_),
    .Y(_12947_));
 sky130_fd_sc_hd__nand2_4 _35512_ (.A(_12595_),
    .B(_12582_),
    .Y(_12948_));
 sky130_fd_sc_hd__a21oi_4 _35513_ (.A1(_12946_),
    .A2(_12947_),
    .B1(_12948_),
    .Y(_12949_));
 sky130_vsdinv _35514_ (.A(_12944_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand2_1 _35515_ (.A(_12940_),
    .B(_12945_),
    .Y(_12951_));
 sky130_fd_sc_hd__o211a_2 _35516_ (.A1(_12950_),
    .A2(_12951_),
    .B1(_12948_),
    .C1(_12946_),
    .X(_12952_));
 sky130_fd_sc_hd__o22ai_4 _35517_ (.A1(_12929_),
    .A2(_12930_),
    .B1(_12949_),
    .B2(_12952_),
    .Y(_12953_));
 sky130_fd_sc_hd__a21oi_4 _35518_ (.A1(_12479_),
    .A2(_12480_),
    .B1(_12559_),
    .Y(_12954_));
 sky130_fd_sc_hd__a21o_1 _35519_ (.A1(_12946_),
    .A2(_12947_),
    .B1(_12948_),
    .X(_12955_));
 sky130_fd_sc_hd__nand3_4 _35520_ (.A(_12946_),
    .B(_12948_),
    .C(_12947_),
    .Y(_12956_));
 sky130_fd_sc_hd__a21o_1 _35521_ (.A1(_12911_),
    .A2(_12917_),
    .B1(_12928_),
    .X(_12957_));
 sky130_fd_sc_hd__nand3_2 _35522_ (.A(_12911_),
    .B(_12917_),
    .C(_12928_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand2_4 _35523_ (.A(_12957_),
    .B(_12958_),
    .Y(_12959_));
 sky130_fd_sc_hd__nand3_4 _35524_ (.A(_12955_),
    .B(_12956_),
    .C(_12959_),
    .Y(_12960_));
 sky130_fd_sc_hd__nand3_4 _35525_ (.A(_12953_),
    .B(_12954_),
    .C(_12960_),
    .Y(_12961_));
 sky130_fd_sc_hd__o21ai_4 _35526_ (.A1(_12593_),
    .A2(_12625_),
    .B1(_12633_),
    .Y(_12962_));
 sky130_fd_sc_hd__and2_1 _35527_ (.A(_12961_),
    .B(_12962_),
    .X(_12963_));
 sky130_fd_sc_hd__nand3b_4 _35528_ (.A_N(_12959_),
    .B(_12955_),
    .C(_12956_),
    .Y(_12964_));
 sky130_fd_sc_hd__o21ai_2 _35529_ (.A1(_12949_),
    .A2(_12952_),
    .B1(_12959_),
    .Y(_12965_));
 sky130_fd_sc_hd__o211ai_4 _35530_ (.A1(_12559_),
    .A2(_12474_),
    .B1(_12964_),
    .C1(_12965_),
    .Y(_12966_));
 sky130_fd_sc_hd__a21oi_4 _35531_ (.A1(_12966_),
    .A2(_12961_),
    .B1(_12962_),
    .Y(_12967_));
 sky130_fd_sc_hd__a21oi_4 _35532_ (.A1(_12963_),
    .A2(_12966_),
    .B1(_12967_),
    .Y(_12968_));
 sky130_fd_sc_hd__nand2_1 _35533_ (.A(_12902_),
    .B(_12968_),
    .Y(_12969_));
 sky130_fd_sc_hd__a21boi_4 _35534_ (.A1(_12647_),
    .A2(_12570_),
    .B1_N(_12563_),
    .Y(_12970_));
 sky130_fd_sc_hd__a22oi_4 _35535_ (.A1(_12470_),
    .A2(_12560_),
    .B1(_12953_),
    .B2(_12960_),
    .Y(_12971_));
 sky130_fd_sc_hd__nand2_1 _35536_ (.A(_12961_),
    .B(_12962_),
    .Y(_12972_));
 sky130_fd_sc_hd__a21o_1 _35537_ (.A1(_12966_),
    .A2(_12961_),
    .B1(_12962_),
    .X(_12973_));
 sky130_fd_sc_hd__o21ai_2 _35538_ (.A1(_12971_),
    .A2(_12972_),
    .B1(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__nand3_2 _35539_ (.A(_12974_),
    .B(_12891_),
    .C(_12901_),
    .Y(_12975_));
 sky130_fd_sc_hd__nand3_4 _35540_ (.A(_12969_),
    .B(_12970_),
    .C(_12975_),
    .Y(_12976_));
 sky130_fd_sc_hd__nand2_1 _35541_ (.A(_12647_),
    .B(_12570_),
    .Y(_12977_));
 sky130_fd_sc_hd__nand2_2 _35542_ (.A(_12977_),
    .B(_12563_),
    .Y(_12978_));
 sky130_fd_sc_hd__nor2_1 _35543_ (.A(_12971_),
    .B(_12972_),
    .Y(_12979_));
 sky130_fd_sc_hd__o2bb2ai_2 _35544_ (.A1_N(_12901_),
    .A2_N(_12891_),
    .B1(_12979_),
    .B2(_12967_),
    .Y(_12980_));
 sky130_fd_sc_hd__nand3_4 _35545_ (.A(_12968_),
    .B(_12891_),
    .C(_12901_),
    .Y(_12981_));
 sky130_fd_sc_hd__nand3_4 _35546_ (.A(_12978_),
    .B(_12980_),
    .C(_12981_),
    .Y(_12982_));
 sky130_vsdinv _35547_ (.A(_12639_),
    .Y(_12983_));
 sky130_fd_sc_hd__nor2_2 _35548_ (.A(_12640_),
    .B(_12635_),
    .Y(_12984_));
 sky130_fd_sc_hd__a22oi_4 _35549_ (.A1(net467),
    .A2(_11587_),
    .B1(_06111_),
    .B2(_11173_),
    .Y(_12985_));
 sky130_fd_sc_hd__nand3_4 _35550_ (.A(_06100_),
    .B(_19915_),
    .C(_20072_),
    .Y(_12986_));
 sky130_fd_sc_hd__nor2_4 _35551_ (.A(_11180_),
    .B(_12986_),
    .Y(_12987_));
 sky130_fd_sc_hd__nand2_2 _35552_ (.A(_05866_),
    .B(\pcpi_mul.rs1[31] ),
    .Y(_12988_));
 sky130_vsdinv _35553_ (.A(_12988_),
    .Y(_12989_));
 sky130_fd_sc_hd__o21ai_2 _35554_ (.A1(_12985_),
    .A2(_12987_),
    .B1(_12989_),
    .Y(_12990_));
 sky130_fd_sc_hd__a22o_1 _35555_ (.A1(_06048_),
    .A2(_09490_),
    .B1(_19906_),
    .B2(_09487_),
    .X(_12991_));
 sky130_fd_sc_hd__a21oi_4 _35556_ (.A1(_12991_),
    .A2(_12615_),
    .B1(_12611_),
    .Y(_12992_));
 sky130_fd_sc_hd__a22o_2 _35557_ (.A1(_05858_),
    .A2(_11587_),
    .B1(_06111_),
    .B2(_20073_),
    .X(_12993_));
 sky130_fd_sc_hd__o211ai_4 _35558_ (.A1(_12688_),
    .A2(_12986_),
    .B1(_12988_),
    .C1(_12993_),
    .Y(_12994_));
 sky130_fd_sc_hd__nand3_4 _35559_ (.A(_12990_),
    .B(_12992_),
    .C(_12994_),
    .Y(_12995_));
 sky130_fd_sc_hd__o21ai_2 _35560_ (.A1(_12985_),
    .A2(_12987_),
    .B1(_12988_),
    .Y(_12996_));
 sky130_fd_sc_hd__o211ai_2 _35561_ (.A1(_12688_),
    .A2(_12986_),
    .B1(_12989_),
    .C1(_12993_),
    .Y(_12997_));
 sky130_fd_sc_hd__nand2_1 _35562_ (.A(_06042_),
    .B(_12102_),
    .Y(_12998_));
 sky130_fd_sc_hd__nand3b_2 _35563_ (.A_N(_12998_),
    .B(_10338_),
    .C(_11927_),
    .Y(_12999_));
 sky130_fd_sc_hd__o21ai_2 _35564_ (.A1(_12613_),
    .A2(_12610_),
    .B1(_12999_),
    .Y(_13000_));
 sky130_fd_sc_hd__nand3_4 _35565_ (.A(_12996_),
    .B(_12997_),
    .C(_13000_),
    .Y(_13001_));
 sky130_fd_sc_hd__nor2_2 _35566_ (.A(_12681_),
    .B(_12679_),
    .Y(_13002_));
 sky130_fd_sc_hd__nor2_4 _35567_ (.A(_12678_),
    .B(_13002_),
    .Y(_13003_));
 sky130_fd_sc_hd__a21oi_2 _35568_ (.A1(_12995_),
    .A2(_13001_),
    .B1(_13003_),
    .Y(_13004_));
 sky130_fd_sc_hd__and3_2 _35569_ (.A(_12995_),
    .B(_13001_),
    .C(_13003_),
    .X(_13005_));
 sky130_fd_sc_hd__a21oi_4 _35570_ (.A1(_12609_),
    .A2(_12617_),
    .B1(_12608_),
    .Y(_13006_));
 sky130_fd_sc_hd__o21ai_4 _35571_ (.A1(_13004_),
    .A2(_13005_),
    .B1(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__o21ai_4 _35572_ (.A1(_12623_),
    .A2(_12620_),
    .B1(_12630_),
    .Y(_13008_));
 sky130_fd_sc_hd__nand3_4 _35573_ (.A(_12995_),
    .B(_13001_),
    .C(_13003_),
    .Y(_13009_));
 sky130_fd_sc_hd__a21o_1 _35574_ (.A1(_12995_),
    .A2(_13001_),
    .B1(_13003_),
    .X(_13010_));
 sky130_fd_sc_hd__nand3_4 _35575_ (.A(_13008_),
    .B(_13009_),
    .C(_13010_),
    .Y(_13011_));
 sky130_fd_sc_hd__a21boi_4 _35576_ (.A1(_12686_),
    .A2(_12694_),
    .B1_N(_12691_),
    .Y(_13012_));
 sky130_vsdinv _35577_ (.A(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__a21o_4 _35578_ (.A1(_13007_),
    .A2(_13011_),
    .B1(_13013_),
    .X(_13014_));
 sky130_fd_sc_hd__nand3_4 _35579_ (.A(_13007_),
    .B(_13011_),
    .C(_13013_),
    .Y(_13015_));
 sky130_vsdinv _35580_ (.A(_12699_),
    .Y(_13016_));
 sky130_fd_sc_hd__o21ai_4 _35581_ (.A1(_13016_),
    .A2(_12697_),
    .B1(_12704_),
    .Y(_13017_));
 sky130_fd_sc_hd__a21o_2 _35582_ (.A1(_13014_),
    .A2(_13015_),
    .B1(_13017_),
    .X(_13018_));
 sky130_fd_sc_hd__nand3_4 _35583_ (.A(_13014_),
    .B(_13017_),
    .C(_13015_),
    .Y(_13019_));
 sky130_fd_sc_hd__a21oi_2 _35584_ (.A1(_12658_),
    .A2(_12660_),
    .B1(_12661_),
    .Y(_13020_));
 sky130_fd_sc_hd__a21o_1 _35585_ (.A1(_12663_),
    .A2(_12355_),
    .B1(_13020_),
    .X(_13021_));
 sky130_fd_sc_hd__nor2_4 _35586_ (.A(net447),
    .B(_19938_),
    .Y(_13022_));
 sky130_fd_sc_hd__a21oi_4 _35587_ (.A1(_19926_),
    .A2(_19938_),
    .B1(_11177_),
    .Y(_13023_));
 sky130_fd_sc_hd__clkinv_8 _35588_ (.A(net503),
    .Y(_13024_));
 sky130_fd_sc_hd__a21oi_2 _35589_ (.A1(_13022_),
    .A2(_12657_),
    .B1(_13024_),
    .Y(_13025_));
 sky130_fd_sc_hd__o31a_1 _35590_ (.A1(_12657_),
    .A2(_13022_),
    .A3(_13023_),
    .B1(_13025_),
    .X(_13026_));
 sky130_fd_sc_hd__nand3_4 _35591_ (.A(_13026_),
    .B(_12351_),
    .C(_12352_),
    .Y(_13027_));
 sky130_vsdinv _35592_ (.A(_13025_),
    .Y(_13028_));
 sky130_fd_sc_hd__nor3_4 _35593_ (.A(_12657_),
    .B(_13022_),
    .C(_13023_),
    .Y(_13029_));
 sky130_fd_sc_hd__o21ai_2 _35594_ (.A1(_13028_),
    .A2(_13029_),
    .B1(_12355_),
    .Y(_13030_));
 sky130_fd_sc_hd__nand2_1 _35595_ (.A(_13027_),
    .B(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__nand2_2 _35596_ (.A(_13021_),
    .B(_13031_),
    .Y(_13032_));
 sky130_fd_sc_hd__a21oi_2 _35597_ (.A1(_12663_),
    .A2(_12355_),
    .B1(_13020_),
    .Y(_13033_));
 sky130_fd_sc_hd__nand3_4 _35598_ (.A(_13033_),
    .B(_13027_),
    .C(_13030_),
    .Y(_13034_));
 sky130_fd_sc_hd__a21o_1 _35599_ (.A1(_13032_),
    .A2(_13034_),
    .B1(_12674_),
    .X(_13035_));
 sky130_fd_sc_hd__nand3_2 _35600_ (.A(_13032_),
    .B(_12674_),
    .C(_13034_),
    .Y(_13036_));
 sky130_fd_sc_hd__nand2_4 _35601_ (.A(_13035_),
    .B(_13036_),
    .Y(_13037_));
 sky130_fd_sc_hd__a21boi_4 _35602_ (.A1(_13018_),
    .A2(_13019_),
    .B1_N(_13037_),
    .Y(_13038_));
 sky130_fd_sc_hd__a21oi_4 _35603_ (.A1(_13014_),
    .A2(_13015_),
    .B1(_13017_),
    .Y(_13039_));
 sky130_fd_sc_hd__and3_1 _35604_ (.A(_13014_),
    .B(_13017_),
    .C(_13015_),
    .X(_13040_));
 sky130_fd_sc_hd__nor3_4 _35605_ (.A(_13037_),
    .B(_13039_),
    .C(_13040_),
    .Y(_13041_));
 sky130_fd_sc_hd__o22ai_4 _35606_ (.A1(_12983_),
    .A2(_12984_),
    .B1(_13038_),
    .B2(_13041_),
    .Y(_13042_));
 sky130_fd_sc_hd__o21ai_2 _35607_ (.A1(_13039_),
    .A2(_13040_),
    .B1(_13037_),
    .Y(_13043_));
 sky130_fd_sc_hd__a31oi_4 _35608_ (.A1(_13014_),
    .A2(_13017_),
    .A3(_13015_),
    .B1(_13037_),
    .Y(_13044_));
 sky130_fd_sc_hd__nand2_4 _35609_ (.A(_13018_),
    .B(_13044_),
    .Y(_13045_));
 sky130_fd_sc_hd__nand2_2 _35610_ (.A(_12641_),
    .B(_12643_),
    .Y(_13046_));
 sky130_fd_sc_hd__nand3_4 _35611_ (.A(_13043_),
    .B(_13045_),
    .C(_13046_),
    .Y(_13047_));
 sky130_fd_sc_hd__nand2_2 _35612_ (.A(_12716_),
    .B(_12715_),
    .Y(_13048_));
 sky130_fd_sc_hd__a21oi_2 _35613_ (.A1(_13042_),
    .A2(_13047_),
    .B1(_13048_),
    .Y(_13049_));
 sky130_fd_sc_hd__and3_1 _35614_ (.A(_13042_),
    .B(_13047_),
    .C(_13048_),
    .X(_13050_));
 sky130_fd_sc_hd__o2bb2ai_4 _35615_ (.A1_N(_12976_),
    .A2_N(_12982_),
    .B1(_13049_),
    .B2(_13050_),
    .Y(_13051_));
 sky130_fd_sc_hd__o2bb2ai_2 _35616_ (.A1_N(_13018_),
    .A2_N(_13044_),
    .B1(_12635_),
    .B2(_12646_),
    .Y(_13052_));
 sky130_fd_sc_hd__nor2_4 _35617_ (.A(_13038_),
    .B(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__nand2_2 _35618_ (.A(_13042_),
    .B(_13048_),
    .Y(_13054_));
 sky130_fd_sc_hd__a21oi_2 _35619_ (.A1(_13043_),
    .A2(_13045_),
    .B1(_13046_),
    .Y(_13055_));
 sky130_fd_sc_hd__o21bai_4 _35620_ (.A1(_13053_),
    .A2(_13055_),
    .B1_N(_13048_),
    .Y(_13056_));
 sky130_fd_sc_hd__o2111ai_4 _35621_ (.A1(_13053_),
    .A2(_13054_),
    .B1(_13056_),
    .C1(_12976_),
    .D1(_12982_),
    .Y(_13057_));
 sky130_vsdinv _35622_ (.A(_12648_),
    .Y(_13058_));
 sky130_fd_sc_hd__nand2_1 _35623_ (.A(_12434_),
    .B(_12645_),
    .Y(_13059_));
 sky130_fd_sc_hd__a21oi_2 _35624_ (.A1(_12645_),
    .A2(_12648_),
    .B1(_12434_),
    .Y(_13060_));
 sky130_fd_sc_hd__nand2_1 _35625_ (.A(_12728_),
    .B(_12722_),
    .Y(_13061_));
 sky130_fd_sc_hd__o22ai_4 _35626_ (.A1(_13058_),
    .A2(_13059_),
    .B1(_13060_),
    .B2(_13061_),
    .Y(_13062_));
 sky130_fd_sc_hd__a21oi_4 _35627_ (.A1(_13051_),
    .A2(_13057_),
    .B1(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__and3_1 _35628_ (.A(_12978_),
    .B(_12980_),
    .C(_12981_),
    .X(_13064_));
 sky130_fd_sc_hd__nand3_2 _35629_ (.A(_13042_),
    .B(_13047_),
    .C(_13048_),
    .Y(_13065_));
 sky130_fd_sc_hd__nand3_4 _35630_ (.A(_12976_),
    .B(_13056_),
    .C(_13065_),
    .Y(_13066_));
 sky130_fd_sc_hd__o211a_2 _35631_ (.A1(_13064_),
    .A2(_13066_),
    .B1(_13051_),
    .C1(_13062_),
    .X(_13067_));
 sky130_vsdinv _35632_ (.A(_12711_),
    .Y(_13068_));
 sky130_fd_sc_hd__nand2_2 _35633_ (.A(_13068_),
    .B(_12671_),
    .Y(_13069_));
 sky130_fd_sc_hd__nand2_2 _35634_ (.A(_12726_),
    .B(_12719_),
    .Y(_13070_));
 sky130_fd_sc_hd__nor2_4 _35635_ (.A(_13069_),
    .B(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__nand2_2 _35636_ (.A(_13070_),
    .B(_13069_),
    .Y(_13072_));
 sky130_vsdinv _35637_ (.A(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__nor2_4 _35638_ (.A(_13071_),
    .B(_13073_),
    .Y(_13074_));
 sky130_fd_sc_hd__o21ai_2 _35639_ (.A1(_13063_),
    .A2(_13067_),
    .B1(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__a22oi_4 _35640_ (.A1(_12742_),
    .A2(_12729_),
    .B1(_12745_),
    .B2(_12752_),
    .Y(_13076_));
 sky130_fd_sc_hd__a21o_2 _35641_ (.A1(_13051_),
    .A2(_13057_),
    .B1(_13062_),
    .X(_13077_));
 sky130_fd_sc_hd__nand3_4 _35642_ (.A(_13062_),
    .B(_13051_),
    .C(_13057_),
    .Y(_13078_));
 sky130_fd_sc_hd__or2b_2 _35643_ (.A(_13071_),
    .B_N(_13072_),
    .X(_13079_));
 sky130_fd_sc_hd__nand3_4 _35644_ (.A(_13077_),
    .B(_13078_),
    .C(_13079_),
    .Y(_13080_));
 sky130_fd_sc_hd__nand3_2 _35645_ (.A(_13075_),
    .B(_13076_),
    .C(_13080_),
    .Y(_13081_));
 sky130_fd_sc_hd__clkbuf_4 _35646_ (.A(_13073_),
    .X(_13082_));
 sky130_fd_sc_hd__o22ai_4 _35647_ (.A1(_13082_),
    .A2(_13071_),
    .B1(_13063_),
    .B2(_13067_),
    .Y(_13083_));
 sky130_fd_sc_hd__nand2_1 _35648_ (.A(_12735_),
    .B(_12724_),
    .Y(_13084_));
 sky130_fd_sc_hd__o22ai_4 _35649_ (.A1(_12739_),
    .A2(_13084_),
    .B1(_12746_),
    .B2(_12736_),
    .Y(_13085_));
 sky130_fd_sc_hd__nand3_2 _35650_ (.A(_13077_),
    .B(_13078_),
    .C(_13074_),
    .Y(_13086_));
 sky130_fd_sc_hd__nand3_4 _35651_ (.A(_13083_),
    .B(_13085_),
    .C(_13086_),
    .Y(_13087_));
 sky130_fd_sc_hd__a21oi_2 _35652_ (.A1(_13081_),
    .A2(_13087_),
    .B1(_12749_),
    .Y(_13088_));
 sky130_fd_sc_hd__and3_1 _35653_ (.A(_13081_),
    .B(_13087_),
    .C(_12749_),
    .X(_13089_));
 sky130_fd_sc_hd__and3_1 _35654_ (.A(_12751_),
    .B(_12753_),
    .C(_12754_),
    .X(_13090_));
 sky130_vsdinv _35655_ (.A(_12405_),
    .Y(_13091_));
 sky130_fd_sc_hd__a31oi_4 _35656_ (.A1(_12425_),
    .A2(_12741_),
    .A3(_12747_),
    .B1(_13091_),
    .Y(_13092_));
 sky130_fd_sc_hd__nor2_2 _35657_ (.A(_13090_),
    .B(_13092_),
    .Y(_13093_));
 sky130_fd_sc_hd__o21ai_4 _35658_ (.A1(_13088_),
    .A2(_13089_),
    .B1(_13093_),
    .Y(_13094_));
 sky130_vsdinv _35659_ (.A(_12749_),
    .Y(_13095_));
 sky130_fd_sc_hd__a31oi_4 _35660_ (.A1(_13075_),
    .A2(_13076_),
    .A3(_13080_),
    .B1(_13095_),
    .Y(_13096_));
 sky130_fd_sc_hd__nand2_1 _35661_ (.A(_13096_),
    .B(_13087_),
    .Y(_13097_));
 sky130_fd_sc_hd__a21o_1 _35662_ (.A1(_13081_),
    .A2(_13087_),
    .B1(_12749_),
    .X(_13098_));
 sky130_fd_sc_hd__o211ai_4 _35663_ (.A1(_13090_),
    .A2(_13092_),
    .B1(_13097_),
    .C1(_13098_),
    .Y(_13099_));
 sky130_fd_sc_hd__nand2_2 _35664_ (.A(_13094_),
    .B(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__nand2_2 _35665_ (.A(_12772_),
    .B(_12764_),
    .Y(_13101_));
 sky130_fd_sc_hd__xnor2_4 _35666_ (.A(_13100_),
    .B(_13101_),
    .Y(_02656_));
 sky130_fd_sc_hd__a21oi_4 _35667_ (.A1(_13077_),
    .A2(_13074_),
    .B1(_13067_),
    .Y(_13102_));
 sky130_fd_sc_hd__nand2_2 _35668_ (.A(_13054_),
    .B(_13047_),
    .Y(_13103_));
 sky130_fd_sc_hd__nand2_1 _35669_ (.A(_13034_),
    .B(_12674_),
    .Y(_13104_));
 sky130_fd_sc_hd__nand2_2 _35670_ (.A(_13104_),
    .B(_13032_),
    .Y(_13105_));
 sky130_vsdinv _35671_ (.A(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__nand2_1 _35672_ (.A(_13103_),
    .B(_13106_),
    .Y(_13107_));
 sky130_vsdinv _35673_ (.A(_13107_),
    .Y(_13108_));
 sky130_fd_sc_hd__nor2_4 _35674_ (.A(_13106_),
    .B(_13103_),
    .Y(_13109_));
 sky130_fd_sc_hd__a21oi_4 _35675_ (.A1(_12888_),
    .A2(_12890_),
    .B1(_12775_),
    .Y(_13110_));
 sky130_fd_sc_hd__o21ai_2 _35676_ (.A1(_12974_),
    .A2(_13110_),
    .B1(_12891_),
    .Y(_13111_));
 sky130_fd_sc_hd__a21oi_2 _35677_ (.A1(_12839_),
    .A2(_12843_),
    .B1(_12836_),
    .Y(_13112_));
 sky130_fd_sc_hd__o21ai_2 _35678_ (.A1(_12899_),
    .A2(_13112_),
    .B1(_12844_),
    .Y(_13113_));
 sky130_fd_sc_hd__a21oi_4 _35679_ (.A1(_12805_),
    .A2(_12809_),
    .B1(_12808_),
    .Y(_13114_));
 sky130_fd_sc_hd__a31oi_4 _35680_ (.A1(_12808_),
    .A2(_12805_),
    .A3(_12809_),
    .B1(_12830_),
    .Y(_13115_));
 sky130_fd_sc_hd__nor2_2 _35681_ (.A(_12791_),
    .B(_12794_),
    .Y(_13116_));
 sky130_fd_sc_hd__nand2_4 _35682_ (.A(_09980_),
    .B(_06696_),
    .Y(_13117_));
 sky130_fd_sc_hd__nand2_4 _35683_ (.A(_09981_),
    .B(_07661_),
    .Y(_13118_));
 sky130_fd_sc_hd__nor2_8 _35684_ (.A(_13117_),
    .B(_13118_),
    .Y(_13119_));
 sky130_fd_sc_hd__nand2_4 _35685_ (.A(_13117_),
    .B(_13118_),
    .Y(_13120_));
 sky130_fd_sc_hd__nand2_2 _35686_ (.A(_08802_),
    .B(_07003_),
    .Y(_13121_));
 sky130_vsdinv _35687_ (.A(_13121_),
    .Y(_13122_));
 sky130_fd_sc_hd__nand3b_4 _35688_ (.A_N(_13119_),
    .B(_13120_),
    .C(_13122_),
    .Y(_13123_));
 sky130_fd_sc_hd__and2_1 _35689_ (.A(_13117_),
    .B(_13118_),
    .X(_13124_));
 sky130_fd_sc_hd__o21ai_2 _35690_ (.A1(_13119_),
    .A2(_13124_),
    .B1(_13121_),
    .Y(_13125_));
 sky130_fd_sc_hd__o211ai_4 _35691_ (.A1(_12790_),
    .A2(_13116_),
    .B1(_13123_),
    .C1(_13125_),
    .Y(_13126_));
 sky130_fd_sc_hd__o21ai_2 _35692_ (.A1(_13119_),
    .A2(_13124_),
    .B1(_13122_),
    .Y(_13127_));
 sky130_fd_sc_hd__nand3b_2 _35693_ (.A_N(_13119_),
    .B(_13120_),
    .C(_13121_),
    .Y(_13128_));
 sky130_fd_sc_hd__a21oi_2 _35694_ (.A1(_12792_),
    .A2(_12795_),
    .B1(_12790_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand3_4 _35695_ (.A(_13127_),
    .B(_13128_),
    .C(_13129_),
    .Y(_13130_));
 sky130_fd_sc_hd__nor2_2 _35696_ (.A(_12814_),
    .B(_12811_),
    .Y(_13131_));
 sky130_fd_sc_hd__nor2_4 _35697_ (.A(_12813_),
    .B(_13131_),
    .Y(_13132_));
 sky130_vsdinv _35698_ (.A(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__a21oi_4 _35699_ (.A1(_13126_),
    .A2(_13130_),
    .B1(_13133_),
    .Y(_13134_));
 sky130_fd_sc_hd__nand2_2 _35700_ (.A(_13126_),
    .B(_13130_),
    .Y(_13135_));
 sky130_fd_sc_hd__nor2_4 _35701_ (.A(_13132_),
    .B(_13135_),
    .Y(_13136_));
 sky130_fd_sc_hd__nor2_4 _35702_ (.A(_13134_),
    .B(_13136_),
    .Y(_13137_));
 sky130_fd_sc_hd__buf_8 _35703_ (.A(_10575_),
    .X(_13138_));
 sky130_fd_sc_hd__buf_6 _35704_ (.A(_18693_),
    .X(_13139_));
 sky130_fd_sc_hd__a22oi_4 _35705_ (.A1(_13138_),
    .A2(_05697_),
    .B1(_05580_),
    .B2(_13139_),
    .Y(_13140_));
 sky130_fd_sc_hd__nand2_8 _35706_ (.A(_19828_),
    .B(_05799_),
    .Y(_13141_));
 sky130_fd_sc_hd__buf_8 _35707_ (.A(_10967_),
    .X(_13142_));
 sky130_fd_sc_hd__nor3_4 _35708_ (.A(_20159_),
    .B(_13141_),
    .C(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__nand2_4 _35709_ (.A(_10573_),
    .B(_05991_),
    .Y(_13144_));
 sky130_vsdinv _35710_ (.A(_13144_),
    .Y(_13145_));
 sky130_fd_sc_hd__o21ai_2 _35711_ (.A1(_13140_),
    .A2(_13143_),
    .B1(_13145_),
    .Y(_13146_));
 sky130_fd_sc_hd__or2b_4 _35712_ (.A(_05474_),
    .B_N(_11778_),
    .X(_13147_));
 sky130_fd_sc_hd__nand2_4 _35713_ (.A(_13147_),
    .B(_13141_),
    .Y(_13148_));
 sky130_fd_sc_hd__nand3b_4 _35714_ (.A_N(_13141_),
    .B(_18694_),
    .C(_05296_),
    .Y(_13149_));
 sky130_fd_sc_hd__nand3_4 _35715_ (.A(_13148_),
    .B(_13149_),
    .C(_13144_),
    .Y(_13150_));
 sky130_fd_sc_hd__a21oi_4 _35716_ (.A1(_12782_),
    .A2(_12780_),
    .B1(_12777_),
    .Y(_13151_));
 sky130_fd_sc_hd__nand3_4 _35717_ (.A(_13146_),
    .B(_13150_),
    .C(_13151_),
    .Y(_13152_));
 sky130_fd_sc_hd__o21ai_2 _35718_ (.A1(_13140_),
    .A2(_13143_),
    .B1(_13144_),
    .Y(_13153_));
 sky130_fd_sc_hd__nand3_4 _35719_ (.A(_13148_),
    .B(_13149_),
    .C(_13145_),
    .Y(_13154_));
 sky130_fd_sc_hd__o21bai_2 _35720_ (.A1(_12779_),
    .A2(_12778_),
    .B1_N(_12777_),
    .Y(_13155_));
 sky130_fd_sc_hd__nand3_4 _35721_ (.A(_13153_),
    .B(_13154_),
    .C(_13155_),
    .Y(_13156_));
 sky130_fd_sc_hd__a22oi_4 _35722_ (.A1(_19836_),
    .A2(net454),
    .B1(_19841_),
    .B2(_20147_),
    .Y(_13157_));
 sky130_fd_sc_hd__nor2_4 _35723_ (.A(_05828_),
    .B(_10983_),
    .Y(_13158_));
 sky130_fd_sc_hd__nand2_2 _35724_ (.A(_09320_),
    .B(_08008_),
    .Y(_13159_));
 sky130_fd_sc_hd__o21ai_2 _35725_ (.A1(_13157_),
    .A2(_13158_),
    .B1(_13159_),
    .Y(_13160_));
 sky130_vsdinv _35726_ (.A(_13160_),
    .Y(_13161_));
 sky130_fd_sc_hd__buf_2 _35727_ (.A(_13158_),
    .X(_13162_));
 sky130_fd_sc_hd__a22o_2 _35728_ (.A1(_19836_),
    .A2(_06148_),
    .B1(_19841_),
    .B2(_10919_),
    .X(_13163_));
 sky130_vsdinv _35729_ (.A(_13159_),
    .Y(_13164_));
 sky130_fd_sc_hd__nand2_2 _35730_ (.A(_13163_),
    .B(_13164_),
    .Y(_13165_));
 sky130_fd_sc_hd__nor2_1 _35731_ (.A(_13162_),
    .B(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__o2bb2ai_2 _35732_ (.A1_N(_13152_),
    .A2_N(_13156_),
    .B1(_13161_),
    .B2(_13166_),
    .Y(_13167_));
 sky130_vsdinv _35733_ (.A(_12787_),
    .Y(_13168_));
 sky130_fd_sc_hd__nand2_1 _35734_ (.A(_12786_),
    .B(_12788_),
    .Y(_13169_));
 sky130_fd_sc_hd__o2bb2ai_2 _35735_ (.A1_N(_12785_),
    .A2_N(_12797_),
    .B1(_13168_),
    .B2(_13169_),
    .Y(_13170_));
 sky130_fd_sc_hd__o21a_1 _35736_ (.A1(_13162_),
    .A2(_13165_),
    .B1(_13160_),
    .X(_13171_));
 sky130_fd_sc_hd__nand3_2 _35737_ (.A(_13152_),
    .B(_13156_),
    .C(_13171_),
    .Y(_13172_));
 sky130_fd_sc_hd__nand3_4 _35738_ (.A(_13167_),
    .B(_13170_),
    .C(_13172_),
    .Y(_13173_));
 sky130_fd_sc_hd__nor2_1 _35739_ (.A(_13157_),
    .B(_13162_),
    .Y(_13174_));
 sky130_fd_sc_hd__nor2_2 _35740_ (.A(_13159_),
    .B(_13174_),
    .Y(_13175_));
 sky130_fd_sc_hd__and2_1 _35741_ (.A(_13174_),
    .B(_13159_),
    .X(_13176_));
 sky130_fd_sc_hd__o2bb2ai_4 _35742_ (.A1_N(_13152_),
    .A2_N(_13156_),
    .B1(_13175_),
    .B2(_13176_),
    .Y(_13177_));
 sky130_fd_sc_hd__a21boi_4 _35743_ (.A1(_12785_),
    .A2(_12797_),
    .B1_N(_12789_),
    .Y(_13178_));
 sky130_fd_sc_hd__o21ai_2 _35744_ (.A1(_13162_),
    .A2(_13165_),
    .B1(_13160_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand3_4 _35745_ (.A(_13152_),
    .B(_13156_),
    .C(_13179_),
    .Y(_13180_));
 sky130_fd_sc_hd__nand3_4 _35746_ (.A(_13177_),
    .B(_13178_),
    .C(_13180_),
    .Y(_13181_));
 sky130_fd_sc_hd__nand3_4 _35747_ (.A(_13137_),
    .B(_13173_),
    .C(_13181_),
    .Y(_13182_));
 sky130_fd_sc_hd__o2bb2ai_2 _35748_ (.A1_N(_13181_),
    .A2_N(_13173_),
    .B1(_13134_),
    .B2(_13136_),
    .Y(_13183_));
 sky130_fd_sc_hd__o211ai_4 _35749_ (.A1(_13114_),
    .A2(_13115_),
    .B1(_13182_),
    .C1(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__nand2_1 _35750_ (.A(_13173_),
    .B(_13181_),
    .Y(_13185_));
 sky130_fd_sc_hd__nand2_1 _35751_ (.A(_13185_),
    .B(_13137_),
    .Y(_13186_));
 sky130_fd_sc_hd__a21oi_4 _35752_ (.A1(_12842_),
    .A2(_12810_),
    .B1(_13114_),
    .Y(_13187_));
 sky130_fd_sc_hd__nand2_1 _35753_ (.A(_13135_),
    .B(_13132_),
    .Y(_13188_));
 sky130_fd_sc_hd__nand3_1 _35754_ (.A(_13126_),
    .B(_13133_),
    .C(_13130_),
    .Y(_13189_));
 sky130_fd_sc_hd__nand2_2 _35755_ (.A(_13188_),
    .B(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__nand3_2 _35756_ (.A(_13173_),
    .B(_13181_),
    .C(_13190_),
    .Y(_13191_));
 sky130_fd_sc_hd__nand3_4 _35757_ (.A(_13186_),
    .B(_13187_),
    .C(_13191_),
    .Y(_13192_));
 sky130_fd_sc_hd__a21oi_4 _35758_ (.A1(_12857_),
    .A2(_12851_),
    .B1(_12849_),
    .Y(_13193_));
 sky130_fd_sc_hd__nand2_2 _35759_ (.A(_08582_),
    .B(_08002_),
    .Y(_13194_));
 sky130_fd_sc_hd__nand2_4 _35760_ (.A(_08577_),
    .B(_06816_),
    .Y(_13195_));
 sky130_fd_sc_hd__nor2_4 _35761_ (.A(_13194_),
    .B(_13195_),
    .Y(_13196_));
 sky130_fd_sc_hd__nand2_2 _35762_ (.A(_13194_),
    .B(_13195_),
    .Y(_13197_));
 sky130_fd_sc_hd__nand2_2 _35763_ (.A(_10435_),
    .B(_07251_),
    .Y(_13198_));
 sky130_vsdinv _35764_ (.A(_13198_),
    .Y(_13199_));
 sky130_fd_sc_hd__nand3b_2 _35765_ (.A_N(_13196_),
    .B(_13197_),
    .C(_13199_),
    .Y(_13200_));
 sky130_fd_sc_hd__and2_1 _35766_ (.A(_13194_),
    .B(_13195_),
    .X(_13201_));
 sky130_fd_sc_hd__o21ai_2 _35767_ (.A1(_13196_),
    .A2(_13201_),
    .B1(_13198_),
    .Y(_13202_));
 sky130_fd_sc_hd__nand3b_4 _35768_ (.A_N(_13193_),
    .B(_13200_),
    .C(_13202_),
    .Y(_13203_));
 sky130_fd_sc_hd__o21ai_2 _35769_ (.A1(_13196_),
    .A2(_13201_),
    .B1(_13199_),
    .Y(_13204_));
 sky130_fd_sc_hd__nand3b_2 _35770_ (.A_N(_13196_),
    .B(_13197_),
    .C(_13198_),
    .Y(_13205_));
 sky130_fd_sc_hd__nand3_4 _35771_ (.A(_13204_),
    .B(_13205_),
    .C(_13193_),
    .Y(_13206_));
 sky130_fd_sc_hd__a22oi_4 _35772_ (.A1(_07483_),
    .A2(_07726_),
    .B1(_19874_),
    .B2(_08060_),
    .Y(_13207_));
 sky130_fd_sc_hd__nand3_4 _35773_ (.A(_12864_),
    .B(_07902_),
    .C(_10113_),
    .Y(_13208_));
 sky130_fd_sc_hd__nor2_4 _35774_ (.A(_10691_),
    .B(_13208_),
    .Y(_13209_));
 sky130_fd_sc_hd__a211o_1 _35775_ (.A1(_19879_),
    .A2(_20112_),
    .B1(_13207_),
    .C1(_13209_),
    .X(_13210_));
 sky130_fd_sc_hd__nand2_2 _35776_ (.A(net457),
    .B(_11492_),
    .Y(_13211_));
 sky130_vsdinv _35777_ (.A(_13211_),
    .Y(_13212_));
 sky130_fd_sc_hd__o21ai_4 _35778_ (.A1(_13207_),
    .A2(_13209_),
    .B1(_13212_),
    .Y(_13213_));
 sky130_fd_sc_hd__nand2_4 _35779_ (.A(_13210_),
    .B(_13213_),
    .Y(_13214_));
 sky130_fd_sc_hd__a21oi_2 _35780_ (.A1(_13203_),
    .A2(_13206_),
    .B1(_13214_),
    .Y(_13215_));
 sky130_fd_sc_hd__nor3_4 _35781_ (.A(_13212_),
    .B(_13207_),
    .C(_13209_),
    .Y(_13216_));
 sky130_vsdinv _35782_ (.A(_13213_),
    .Y(_13217_));
 sky130_fd_sc_hd__o211a_2 _35783_ (.A1(_13216_),
    .A2(_13217_),
    .B1(_13206_),
    .C1(_13203_),
    .X(_13218_));
 sky130_fd_sc_hd__nand2_4 _35784_ (.A(_12841_),
    .B(_12825_),
    .Y(_13219_));
 sky130_fd_sc_hd__o21bai_4 _35785_ (.A1(_13215_),
    .A2(_13218_),
    .B1_N(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__a21o_1 _35786_ (.A1(_13203_),
    .A2(_13206_),
    .B1(_13214_),
    .X(_13221_));
 sky130_fd_sc_hd__nand3_4 _35787_ (.A(_13203_),
    .B(_13214_),
    .C(_13206_),
    .Y(_13222_));
 sky130_fd_sc_hd__nand3_4 _35788_ (.A(_13221_),
    .B(_13219_),
    .C(_13222_),
    .Y(_13223_));
 sky130_fd_sc_hd__nand2_2 _35789_ (.A(_12880_),
    .B(_12863_),
    .Y(_13224_));
 sky130_fd_sc_hd__a21oi_4 _35790_ (.A1(_13220_),
    .A2(_13223_),
    .B1(_13224_),
    .Y(_13225_));
 sky130_fd_sc_hd__nand3_2 _35791_ (.A(_13220_),
    .B(_13223_),
    .C(_13224_),
    .Y(_13226_));
 sky130_vsdinv _35792_ (.A(_13226_),
    .Y(_13227_));
 sky130_fd_sc_hd__o2bb2ai_1 _35793_ (.A1_N(_13184_),
    .A2_N(_13192_),
    .B1(_13225_),
    .B2(_13227_),
    .Y(_13228_));
 sky130_vsdinv _35794_ (.A(_13224_),
    .Y(_13229_));
 sky130_fd_sc_hd__a21oi_4 _35795_ (.A1(_13221_),
    .A2(_13222_),
    .B1(_13219_),
    .Y(_13230_));
 sky130_fd_sc_hd__nor2_2 _35796_ (.A(_13229_),
    .B(_13230_),
    .Y(_13231_));
 sky130_fd_sc_hd__a21oi_4 _35797_ (.A1(_13231_),
    .A2(_13223_),
    .B1(_13225_),
    .Y(_13232_));
 sky130_fd_sc_hd__nand3_2 _35798_ (.A(_13232_),
    .B(_13192_),
    .C(_13184_),
    .Y(_13233_));
 sky130_fd_sc_hd__nand3_4 _35799_ (.A(_13113_),
    .B(_13228_),
    .C(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__nand2_1 _35800_ (.A(_13192_),
    .B(_13184_),
    .Y(_13235_));
 sky130_fd_sc_hd__nand2_1 _35801_ (.A(_13235_),
    .B(_13232_),
    .Y(_13236_));
 sky130_fd_sc_hd__a21boi_2 _35802_ (.A1(_12889_),
    .A2(_12834_),
    .B1_N(_12844_),
    .Y(_13237_));
 sky130_fd_sc_hd__a21o_1 _35803_ (.A1(_13220_),
    .A2(_13223_),
    .B1(_13224_),
    .X(_13238_));
 sky130_fd_sc_hd__nand2_2 _35804_ (.A(_13238_),
    .B(_13226_),
    .Y(_13239_));
 sky130_fd_sc_hd__nand3_2 _35805_ (.A(_13239_),
    .B(_13192_),
    .C(_13184_),
    .Y(_13240_));
 sky130_fd_sc_hd__nand3_4 _35806_ (.A(_13236_),
    .B(_13237_),
    .C(_13240_),
    .Y(_13241_));
 sky130_fd_sc_hd__a31o_2 _35807_ (.A1(_12941_),
    .A2(_12943_),
    .A3(_12942_),
    .B1(_12945_),
    .X(_13242_));
 sky130_fd_sc_hd__o21ba_2 _35808_ (.A1(_12865_),
    .A2(_12868_),
    .B1_N(_12866_),
    .X(_13243_));
 sky130_fd_sc_hd__nand2_2 _35809_ (.A(_11092_),
    .B(_08453_),
    .Y(_13244_));
 sky130_fd_sc_hd__nand2_4 _35810_ (.A(_12576_),
    .B(_09926_),
    .Y(_13245_));
 sky130_fd_sc_hd__or2_2 _35811_ (.A(_13244_),
    .B(_13245_),
    .X(_13246_));
 sky130_fd_sc_hd__nand2_2 _35812_ (.A(_13244_),
    .B(_13245_),
    .Y(_13247_));
 sky130_fd_sc_hd__nand2_2 _35813_ (.A(_06641_),
    .B(_10811_),
    .Y(_13248_));
 sky130_fd_sc_hd__nand3_4 _35814_ (.A(_13246_),
    .B(_13247_),
    .C(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__nor2_4 _35815_ (.A(_13244_),
    .B(_13245_),
    .Y(_13250_));
 sky130_fd_sc_hd__and2_2 _35816_ (.A(_13244_),
    .B(_13245_),
    .X(_13251_));
 sky130_vsdinv _35817_ (.A(_13248_),
    .Y(_13252_));
 sky130_fd_sc_hd__o21ai_2 _35818_ (.A1(_13250_),
    .A2(_13251_),
    .B1(_13252_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand3_1 _35819_ (.A(_13243_),
    .B(_13249_),
    .C(_13253_),
    .Y(_13254_));
 sky130_fd_sc_hd__o21ai_2 _35820_ (.A1(_13250_),
    .A2(_13251_),
    .B1(_13248_),
    .Y(_13255_));
 sky130_fd_sc_hd__nand3_4 _35821_ (.A(_13246_),
    .B(_13247_),
    .C(_13252_),
    .Y(_13256_));
 sky130_fd_sc_hd__o21bai_4 _35822_ (.A1(_12865_),
    .A2(_12868_),
    .B1_N(_12866_),
    .Y(_13257_));
 sky130_fd_sc_hd__nand3_4 _35823_ (.A(_13255_),
    .B(_13256_),
    .C(_13257_),
    .Y(_13258_));
 sky130_fd_sc_hd__a21oi_4 _35824_ (.A1(_12938_),
    .A2(_12935_),
    .B1(_12933_),
    .Y(_13259_));
 sky130_vsdinv _35825_ (.A(_13259_),
    .Y(_13260_));
 sky130_fd_sc_hd__a21o_2 _35826_ (.A1(_13254_),
    .A2(_13258_),
    .B1(_13260_),
    .X(_13261_));
 sky130_fd_sc_hd__a31oi_4 _35827_ (.A1(_13243_),
    .A2(_13253_),
    .A3(_13249_),
    .B1(_13259_),
    .Y(_13262_));
 sky130_fd_sc_hd__nand2_4 _35828_ (.A(_13262_),
    .B(_13258_),
    .Y(_13263_));
 sky130_fd_sc_hd__a22oi_4 _35829_ (.A1(_12940_),
    .A2(_13242_),
    .B1(_13261_),
    .B2(_13263_),
    .Y(_13264_));
 sky130_vsdinv _35830_ (.A(_12951_),
    .Y(_13265_));
 sky130_fd_sc_hd__o211a_1 _35831_ (.A1(_12950_),
    .A2(_13265_),
    .B1(_13263_),
    .C1(_13261_),
    .X(_13266_));
 sky130_fd_sc_hd__nand2_4 _35832_ (.A(_11058_),
    .B(_09041_),
    .Y(_13267_));
 sky130_fd_sc_hd__nand2_4 _35833_ (.A(_07422_),
    .B(_09038_),
    .Y(_13268_));
 sky130_fd_sc_hd__nor2_8 _35834_ (.A(_13267_),
    .B(_13268_),
    .Y(_13269_));
 sky130_fd_sc_hd__and2_1 _35835_ (.A(_13267_),
    .B(_13268_),
    .X(_13270_));
 sky130_fd_sc_hd__clkinv_8 _35836_ (.A(net505),
    .Y(_13271_));
 sky130_fd_sc_hd__nor2_4 _35837_ (.A(_13271_),
    .B(_10780_),
    .Y(_13272_));
 sky130_fd_sc_hd__o21bai_4 _35838_ (.A1(_13269_),
    .A2(_13270_),
    .B1_N(_13272_),
    .Y(_13273_));
 sky130_fd_sc_hd__nand2_2 _35839_ (.A(_12907_),
    .B(_12915_),
    .Y(_13274_));
 sky130_fd_sc_hd__nand2_4 _35840_ (.A(_13267_),
    .B(_13268_),
    .Y(_13275_));
 sky130_fd_sc_hd__nand3b_4 _35841_ (.A_N(_13269_),
    .B(_13272_),
    .C(_13275_),
    .Y(_13276_));
 sky130_fd_sc_hd__nand3_4 _35842_ (.A(_13273_),
    .B(_13274_),
    .C(_13276_),
    .Y(_13277_));
 sky130_vsdinv _35843_ (.A(_13277_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand2_1 _35844_ (.A(_13273_),
    .B(_13276_),
    .Y(_13279_));
 sky130_fd_sc_hd__a22oi_4 _35845_ (.A1(_19903_),
    .A2(_20087_),
    .B1(_19907_),
    .B2(_11165_),
    .Y(_13280_));
 sky130_fd_sc_hd__nand2_2 _35846_ (.A(_06119_),
    .B(_09787_),
    .Y(_13281_));
 sky130_fd_sc_hd__nand2_2 _35847_ (.A(_10347_),
    .B(_11157_),
    .Y(_13282_));
 sky130_fd_sc_hd__nor2_4 _35848_ (.A(_13281_),
    .B(_13282_),
    .Y(_13283_));
 sky130_fd_sc_hd__nor2_1 _35849_ (.A(_13280_),
    .B(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__nor2_2 _35850_ (.A(_05633_),
    .B(_12688_),
    .Y(_13285_));
 sky130_fd_sc_hd__nand2_1 _35851_ (.A(_13284_),
    .B(_13285_),
    .Y(_13286_));
 sky130_fd_sc_hd__o21bai_2 _35852_ (.A1(_13280_),
    .A2(_13283_),
    .B1_N(_13285_),
    .Y(_13287_));
 sky130_fd_sc_hd__nand2_4 _35853_ (.A(_13286_),
    .B(_13287_),
    .Y(_13288_));
 sky130_fd_sc_hd__a31o_1 _35854_ (.A1(_13279_),
    .A2(_12915_),
    .A3(_12907_),
    .B1(_13288_),
    .X(_13289_));
 sky130_fd_sc_hd__a21oi_4 _35855_ (.A1(_13273_),
    .A2(_13276_),
    .B1(_13274_),
    .Y(_13290_));
 sky130_fd_sc_hd__o21ai_2 _35856_ (.A1(_13290_),
    .A2(_13278_),
    .B1(_13288_),
    .Y(_13291_));
 sky130_fd_sc_hd__o21a_2 _35857_ (.A1(_13278_),
    .A2(_13289_),
    .B1(_13291_),
    .X(_13292_));
 sky130_fd_sc_hd__o21ai_4 _35858_ (.A1(_13264_),
    .A2(_13266_),
    .B1(_13292_),
    .Y(_13293_));
 sky130_fd_sc_hd__a21boi_4 _35859_ (.A1(_12877_),
    .A2(_12884_),
    .B1_N(_12882_),
    .Y(_13294_));
 sky130_fd_sc_hd__a22o_2 _35860_ (.A1(_12940_),
    .A2(_13242_),
    .B1(_13261_),
    .B2(_13263_),
    .X(_13295_));
 sky130_fd_sc_hd__o21ai_4 _35861_ (.A1(_13278_),
    .A2(_13289_),
    .B1(_13291_),
    .Y(_13296_));
 sky130_fd_sc_hd__o211ai_4 _35862_ (.A1(_12950_),
    .A2(_13265_),
    .B1(_13263_),
    .C1(_13261_),
    .Y(_13297_));
 sky130_fd_sc_hd__nand3_4 _35863_ (.A(_13295_),
    .B(_13296_),
    .C(_13297_),
    .Y(_13298_));
 sky130_fd_sc_hd__nand3_4 _35864_ (.A(_13293_),
    .B(_13294_),
    .C(_13298_),
    .Y(_13299_));
 sky130_fd_sc_hd__o21ai_2 _35865_ (.A1(_13264_),
    .A2(_13266_),
    .B1(_13296_),
    .Y(_13300_));
 sky130_fd_sc_hd__nand2_2 _35866_ (.A(_12898_),
    .B(_12882_),
    .Y(_13301_));
 sky130_fd_sc_hd__nand3_4 _35867_ (.A(_13295_),
    .B(_13292_),
    .C(_13297_),
    .Y(_13302_));
 sky130_fd_sc_hd__nand3_4 _35868_ (.A(_13300_),
    .B(_13301_),
    .C(_13302_),
    .Y(_13303_));
 sky130_fd_sc_hd__nor2_2 _35869_ (.A(_12959_),
    .B(_12949_),
    .Y(_13304_));
 sky130_fd_sc_hd__or2_4 _35870_ (.A(_12952_),
    .B(_13304_),
    .X(_13305_));
 sky130_fd_sc_hd__a21oi_4 _35871_ (.A1(_13299_),
    .A2(_13303_),
    .B1(_13305_),
    .Y(_13306_));
 sky130_fd_sc_hd__and3_1 _35872_ (.A(_13299_),
    .B(_13303_),
    .C(_13305_),
    .X(_13307_));
 sky130_fd_sc_hd__o2bb2ai_2 _35873_ (.A1_N(_13234_),
    .A2_N(_13241_),
    .B1(_13306_),
    .B2(_13307_),
    .Y(_13308_));
 sky130_fd_sc_hd__o2bb2ai_1 _35874_ (.A1_N(_13299_),
    .A2_N(_13303_),
    .B1(_12952_),
    .B2(_13304_),
    .Y(_13309_));
 sky130_fd_sc_hd__nor2_2 _35875_ (.A(_12952_),
    .B(_13304_),
    .Y(_13310_));
 sky130_fd_sc_hd__nand3_1 _35876_ (.A(_13299_),
    .B(_13303_),
    .C(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__nand2_2 _35877_ (.A(_13309_),
    .B(_13311_),
    .Y(_13312_));
 sky130_fd_sc_hd__nand3_4 _35878_ (.A(_13312_),
    .B(_13234_),
    .C(_13241_),
    .Y(_13313_));
 sky130_fd_sc_hd__nand3_4 _35879_ (.A(_13111_),
    .B(_13308_),
    .C(_13313_),
    .Y(_13314_));
 sky130_fd_sc_hd__nand2_1 _35880_ (.A(_13241_),
    .B(_13234_),
    .Y(_13315_));
 sky130_fd_sc_hd__nand2_1 _35881_ (.A(_13315_),
    .B(_13312_),
    .Y(_13316_));
 sky130_fd_sc_hd__a21boi_4 _35882_ (.A1(_12968_),
    .A2(_12901_),
    .B1_N(_12891_),
    .Y(_13317_));
 sky130_fd_sc_hd__o211ai_4 _35883_ (.A1(_13306_),
    .A2(_13307_),
    .B1(_13234_),
    .C1(_13241_),
    .Y(_13318_));
 sky130_fd_sc_hd__nand3_4 _35884_ (.A(_13316_),
    .B(_13317_),
    .C(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__a22oi_4 _35885_ (.A1(_06096_),
    .A2(_10760_),
    .B1(_06098_),
    .B2(_20069_),
    .Y(_13320_));
 sky130_fd_sc_hd__nand3_4 _35886_ (.A(_19912_),
    .B(_06474_),
    .C(_10777_),
    .Y(_13321_));
 sky130_fd_sc_hd__nor2_4 _35887_ (.A(_10772_),
    .B(_13321_),
    .Y(_13322_));
 sky130_fd_sc_hd__nand2_2 _35888_ (.A(\pcpi_mul.rs1[32] ),
    .B(_05865_),
    .Y(_13323_));
 sky130_vsdinv _35889_ (.A(_13323_),
    .Y(_13324_));
 sky130_fd_sc_hd__clkbuf_4 _35890_ (.A(_13324_),
    .X(_13325_));
 sky130_fd_sc_hd__o21ai_2 _35891_ (.A1(_13320_),
    .A2(_13322_),
    .B1(_13325_),
    .Y(_13326_));
 sky130_fd_sc_hd__o21ai_1 _35892_ (.A1(_12920_),
    .A2(_12921_),
    .B1(_12923_),
    .Y(_13327_));
 sky130_fd_sc_hd__nand2_1 _35893_ (.A(_13327_),
    .B(_12926_),
    .Y(_13328_));
 sky130_fd_sc_hd__buf_4 _35894_ (.A(_13323_),
    .X(_13329_));
 sky130_fd_sc_hd__a22o_1 _35895_ (.A1(_10809_),
    .A2(_10760_),
    .B1(_11206_),
    .B2(_20069_),
    .X(_13330_));
 sky130_fd_sc_hd__o211ai_2 _35896_ (.A1(_10767_),
    .A2(_13321_),
    .B1(_13329_),
    .C1(_13330_),
    .Y(_13331_));
 sky130_fd_sc_hd__nand3_4 _35897_ (.A(_13326_),
    .B(_13328_),
    .C(_13331_),
    .Y(_13332_));
 sky130_fd_sc_hd__o21ai_2 _35898_ (.A1(_13320_),
    .A2(_13322_),
    .B1(_13329_),
    .Y(_13333_));
 sky130_fd_sc_hd__o21ai_2 _35899_ (.A1(_12923_),
    .A2(_12919_),
    .B1(_12925_),
    .Y(_13334_));
 sky130_fd_sc_hd__o211ai_2 _35900_ (.A1(_10767_),
    .A2(_13321_),
    .B1(_13325_),
    .C1(_13330_),
    .Y(_13335_));
 sky130_fd_sc_hd__nand3_4 _35901_ (.A(_13333_),
    .B(_13334_),
    .C(_13335_),
    .Y(_13336_));
 sky130_fd_sc_hd__nor2_4 _35902_ (.A(_12989_),
    .B(_12987_),
    .Y(_13337_));
 sky130_fd_sc_hd__o2bb2ai_4 _35903_ (.A1_N(_13332_),
    .A2_N(_13336_),
    .B1(_12985_),
    .B2(_13337_),
    .Y(_13338_));
 sky130_fd_sc_hd__nor2_2 _35904_ (.A(_12985_),
    .B(_13337_),
    .Y(_13339_));
 sky130_fd_sc_hd__nand3_4 _35905_ (.A(_13332_),
    .B(_13336_),
    .C(_13339_),
    .Y(_13340_));
 sky130_fd_sc_hd__nand2_1 _35906_ (.A(_12917_),
    .B(_12928_),
    .Y(_13341_));
 sky130_fd_sc_hd__nand2_4 _35907_ (.A(_13341_),
    .B(_12911_),
    .Y(_13342_));
 sky130_fd_sc_hd__a21oi_4 _35908_ (.A1(_13338_),
    .A2(_13340_),
    .B1(_13342_),
    .Y(_13343_));
 sky130_vsdinv _35909_ (.A(_13336_),
    .Y(_13344_));
 sky130_fd_sc_hd__nand2_1 _35910_ (.A(_13332_),
    .B(_13339_),
    .Y(_13345_));
 sky130_fd_sc_hd__o211a_1 _35911_ (.A1(_13344_),
    .A2(_13345_),
    .B1(_13338_),
    .C1(_13342_),
    .X(_13346_));
 sky130_fd_sc_hd__nand2_1 _35912_ (.A(_12995_),
    .B(_13003_),
    .Y(_13347_));
 sky130_fd_sc_hd__nand2_2 _35913_ (.A(_13347_),
    .B(_13001_),
    .Y(_13348_));
 sky130_fd_sc_hd__o21ai_2 _35914_ (.A1(_13343_),
    .A2(_13346_),
    .B1(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__a21boi_2 _35915_ (.A1(_13007_),
    .A2(_13013_),
    .B1_N(_13011_),
    .Y(_13350_));
 sky130_fd_sc_hd__a21o_1 _35916_ (.A1(_13338_),
    .A2(_13340_),
    .B1(_13342_),
    .X(_13351_));
 sky130_fd_sc_hd__nand3_4 _35917_ (.A(_13342_),
    .B(_13338_),
    .C(_13340_),
    .Y(_13352_));
 sky130_vsdinv _35918_ (.A(_13348_),
    .Y(_13353_));
 sky130_fd_sc_hd__nand3_2 _35919_ (.A(_13351_),
    .B(_13352_),
    .C(_13353_),
    .Y(_13354_));
 sky130_fd_sc_hd__nand3_4 _35920_ (.A(_13349_),
    .B(_13350_),
    .C(_13354_),
    .Y(_13355_));
 sky130_fd_sc_hd__o21ai_2 _35921_ (.A1(_13343_),
    .A2(_13346_),
    .B1(_13353_),
    .Y(_13356_));
 sky130_fd_sc_hd__nand2_1 _35922_ (.A(_13008_),
    .B(_13010_),
    .Y(_13357_));
 sky130_fd_sc_hd__a21oi_2 _35923_ (.A1(_13010_),
    .A2(_13009_),
    .B1(_13008_),
    .Y(_13358_));
 sky130_fd_sc_hd__o22ai_4 _35924_ (.A1(_13005_),
    .A2(_13357_),
    .B1(_13012_),
    .B2(_13358_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand3_2 _35925_ (.A(_13351_),
    .B(_13352_),
    .C(_13348_),
    .Y(_13360_));
 sky130_fd_sc_hd__nand3_4 _35926_ (.A(_13356_),
    .B(_13359_),
    .C(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand2_1 _35927_ (.A(_13355_),
    .B(_13361_),
    .Y(_13362_));
 sky130_vsdinv _35928_ (.A(_13030_),
    .Y(_13363_));
 sky130_fd_sc_hd__nor2_1 _35929_ (.A(_13028_),
    .B(_13363_),
    .Y(_13364_));
 sky130_fd_sc_hd__a21o_1 _35930_ (.A1(_12356_),
    .A2(_13028_),
    .B1(_12673_),
    .X(_13365_));
 sky130_fd_sc_hd__nand2_1 _35931_ (.A(_13363_),
    .B(_13025_),
    .Y(_13366_));
 sky130_fd_sc_hd__nand2_2 _35932_ (.A(_12353_),
    .B(_13028_),
    .Y(_13367_));
 sky130_fd_sc_hd__nand3_2 _35933_ (.A(_13366_),
    .B(_12674_),
    .C(_13367_),
    .Y(_13368_));
 sky130_fd_sc_hd__o21a_1 _35934_ (.A1(_13364_),
    .A2(_13365_),
    .B1(_13368_),
    .X(_13369_));
 sky130_vsdinv _35935_ (.A(_13369_),
    .Y(_13370_));
 sky130_fd_sc_hd__nand2_1 _35936_ (.A(_13362_),
    .B(_13370_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand2_1 _35937_ (.A(_12972_),
    .B(_12966_),
    .Y(_13372_));
 sky130_fd_sc_hd__nand3_2 _35938_ (.A(_13355_),
    .B(_13361_),
    .C(_13369_),
    .Y(_13373_));
 sky130_fd_sc_hd__nand3_4 _35939_ (.A(_13371_),
    .B(_13372_),
    .C(_13373_),
    .Y(_13374_));
 sky130_fd_sc_hd__buf_2 _35940_ (.A(_13374_),
    .X(_13375_));
 sky130_fd_sc_hd__nand2_1 _35941_ (.A(_13362_),
    .B(_13369_),
    .Y(_13376_));
 sky130_fd_sc_hd__a21oi_2 _35942_ (.A1(_12961_),
    .A2(_12962_),
    .B1(_12971_),
    .Y(_13377_));
 sky130_fd_sc_hd__nand3_2 _35943_ (.A(_13355_),
    .B(_13370_),
    .C(_13361_),
    .Y(_13378_));
 sky130_fd_sc_hd__nand3_4 _35944_ (.A(_13376_),
    .B(_13377_),
    .C(_13378_),
    .Y(_13379_));
 sky130_fd_sc_hd__nand2_4 _35945_ (.A(_13045_),
    .B(_13019_),
    .Y(_13380_));
 sky130_fd_sc_hd__a21oi_4 _35946_ (.A1(_13375_),
    .A2(_13379_),
    .B1(_13380_),
    .Y(_13381_));
 sky130_fd_sc_hd__nand3_4 _35947_ (.A(_13374_),
    .B(_13379_),
    .C(_13380_),
    .Y(_13382_));
 sky130_vsdinv _35948_ (.A(_13382_),
    .Y(_13383_));
 sky130_fd_sc_hd__o2bb2ai_4 _35949_ (.A1_N(_13314_),
    .A2_N(_13319_),
    .B1(_13381_),
    .B2(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__and2_1 _35950_ (.A(_13379_),
    .B(_13380_),
    .X(_13385_));
 sky130_fd_sc_hd__a21oi_4 _35951_ (.A1(_13385_),
    .A2(_13375_),
    .B1(_13381_),
    .Y(_13386_));
 sky130_fd_sc_hd__nand3_4 _35952_ (.A(_13386_),
    .B(_13314_),
    .C(_13319_),
    .Y(_13387_));
 sky130_fd_sc_hd__nand2_4 _35953_ (.A(_13066_),
    .B(_12982_),
    .Y(_13388_));
 sky130_fd_sc_hd__a21oi_4 _35954_ (.A1(_13384_),
    .A2(_13387_),
    .B1(_13388_),
    .Y(_13389_));
 sky130_fd_sc_hd__nand2_1 _35955_ (.A(_13308_),
    .B(_13313_),
    .Y(_13390_));
 sky130_fd_sc_hd__nand2_1 _35956_ (.A(_13375_),
    .B(_13379_),
    .Y(_13391_));
 sky130_fd_sc_hd__nor2_1 _35957_ (.A(_13040_),
    .B(_13041_),
    .Y(_13392_));
 sky130_fd_sc_hd__nand2_1 _35958_ (.A(_13391_),
    .B(_13392_),
    .Y(_13393_));
 sky130_fd_sc_hd__nand2_1 _35959_ (.A(_13393_),
    .B(_13382_),
    .Y(_13394_));
 sky130_fd_sc_hd__a21oi_1 _35960_ (.A1(_13390_),
    .A2(_13317_),
    .B1(_13394_),
    .Y(_13395_));
 sky130_fd_sc_hd__a2bb2oi_1 _35961_ (.A1_N(_13381_),
    .A2_N(_13383_),
    .B1(_13314_),
    .B2(_13319_),
    .Y(_13396_));
 sky130_fd_sc_hd__a221oi_2 _35962_ (.A1(_13066_),
    .A2(_12982_),
    .B1(_13395_),
    .B2(_13314_),
    .C1(_13396_),
    .Y(_13397_));
 sky130_fd_sc_hd__o22ai_4 _35963_ (.A1(_13108_),
    .A2(_13109_),
    .B1(_13389_),
    .B2(_13397_),
    .Y(_13398_));
 sky130_fd_sc_hd__a21o_1 _35964_ (.A1(_13384_),
    .A2(_13387_),
    .B1(_13388_),
    .X(_13399_));
 sky130_fd_sc_hd__nand3_4 _35965_ (.A(_13388_),
    .B(_13384_),
    .C(_13387_),
    .Y(_13400_));
 sky130_fd_sc_hd__and2b_2 _35966_ (.A_N(_13109_),
    .B(_13107_),
    .X(_13401_));
 sky130_fd_sc_hd__nand3_4 _35967_ (.A(_13399_),
    .B(_13400_),
    .C(_13401_),
    .Y(_13402_));
 sky130_fd_sc_hd__nand3_4 _35968_ (.A(_13102_),
    .B(_13398_),
    .C(_13402_),
    .Y(_13403_));
 sky130_vsdinv _35969_ (.A(_13103_),
    .Y(_13404_));
 sky130_fd_sc_hd__nor2_8 _35970_ (.A(_13106_),
    .B(_13404_),
    .Y(_13405_));
 sky130_fd_sc_hd__nor2_2 _35971_ (.A(_13105_),
    .B(_13103_),
    .Y(_13406_));
 sky130_fd_sc_hd__o22ai_4 _35972_ (.A1(_13405_),
    .A2(_13406_),
    .B1(_13389_),
    .B2(_13397_),
    .Y(_13407_));
 sky130_fd_sc_hd__o211ai_4 _35973_ (.A1(_13108_),
    .A2(_13109_),
    .B1(_13400_),
    .C1(_13399_),
    .Y(_13408_));
 sky130_fd_sc_hd__o21ai_2 _35974_ (.A1(_13079_),
    .A2(_13063_),
    .B1(_13078_),
    .Y(_13409_));
 sky130_fd_sc_hd__nand3_4 _35975_ (.A(_13407_),
    .B(_13408_),
    .C(_13409_),
    .Y(_13410_));
 sky130_fd_sc_hd__a21oi_2 _35976_ (.A1(_13403_),
    .A2(_13410_),
    .B1(_13082_),
    .Y(_13411_));
 sky130_fd_sc_hd__and3_1 _35977_ (.A(_13403_),
    .B(_13410_),
    .C(_13082_),
    .X(_13412_));
 sky130_vsdinv _35978_ (.A(_13087_),
    .Y(_13413_));
 sky130_fd_sc_hd__nor2_2 _35979_ (.A(_13096_),
    .B(_13413_),
    .Y(_13414_));
 sky130_fd_sc_hd__o21ai_4 _35980_ (.A1(_13411_),
    .A2(_13412_),
    .B1(_13414_),
    .Y(_13415_));
 sky130_fd_sc_hd__nand3_4 _35981_ (.A(_13403_),
    .B(_13410_),
    .C(_13082_),
    .Y(_13416_));
 sky130_fd_sc_hd__a21o_1 _35982_ (.A1(_13403_),
    .A2(_13410_),
    .B1(_13082_),
    .X(_13417_));
 sky130_fd_sc_hd__o211ai_4 _35983_ (.A1(_13413_),
    .A2(_13096_),
    .B1(_13416_),
    .C1(_13417_),
    .Y(_13418_));
 sky130_fd_sc_hd__nand2_2 _35984_ (.A(_13415_),
    .B(_13418_),
    .Y(_13419_));
 sky130_fd_sc_hd__nand2_1 _35985_ (.A(_12760_),
    .B(_12763_),
    .Y(_13420_));
 sky130_fd_sc_hd__o2111ai_4 _35986_ (.A1(_12756_),
    .A2(_13420_),
    .B1(_13099_),
    .C1(_13094_),
    .D1(_12761_),
    .Y(_13421_));
 sky130_fd_sc_hd__nand2_1 _35987_ (.A(_12764_),
    .B(_13099_),
    .Y(_13422_));
 sky130_fd_sc_hd__nand2_2 _35988_ (.A(_13422_),
    .B(_13094_),
    .Y(_13423_));
 sky130_fd_sc_hd__o21ai_4 _35989_ (.A1(_13421_),
    .A2(_12771_),
    .B1(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__xnor2_4 _35990_ (.A(_13419_),
    .B(_13424_),
    .Y(_02657_));
 sky130_fd_sc_hd__and3_1 _35991_ (.A(_13255_),
    .B(_13256_),
    .C(_13257_),
    .X(_13425_));
 sky130_fd_sc_hd__and4_2 _35992_ (.A(_11092_),
    .B(_19887_),
    .C(_08881_),
    .D(_08884_),
    .X(_13426_));
 sky130_fd_sc_hd__a22o_1 _35993_ (.A1(_19882_),
    .A2(_11078_),
    .B1(_11455_),
    .B2(_20102_),
    .X(_13427_));
 sky130_fd_sc_hd__nand2_2 _35994_ (.A(_06641_),
    .B(_11503_),
    .Y(_13428_));
 sky130_fd_sc_hd__nand3b_2 _35995_ (.A_N(_13426_),
    .B(_13427_),
    .C(_13428_),
    .Y(_13429_));
 sky130_fd_sc_hd__o22a_1 _35996_ (.A1(_10704_),
    .A2(_13208_),
    .B1(_13211_),
    .B2(_13207_),
    .X(_13430_));
 sky130_fd_sc_hd__a22oi_4 _35997_ (.A1(_19882_),
    .A2(_11078_),
    .B1(_19888_),
    .B2(_12303_),
    .Y(_13431_));
 sky130_vsdinv _35998_ (.A(_13428_),
    .Y(_13432_));
 sky130_fd_sc_hd__o21ai_2 _35999_ (.A1(_13431_),
    .A2(_13426_),
    .B1(_13432_),
    .Y(_13433_));
 sky130_fd_sc_hd__nand3_4 _36000_ (.A(_13429_),
    .B(_13430_),
    .C(_13433_),
    .Y(_13434_));
 sky130_fd_sc_hd__nand3b_2 _36001_ (.A_N(_13426_),
    .B(_13427_),
    .C(_13432_),
    .Y(_13435_));
 sky130_fd_sc_hd__o22ai_4 _36002_ (.A1(_10704_),
    .A2(_13208_),
    .B1(_13211_),
    .B2(_13207_),
    .Y(_13436_));
 sky130_fd_sc_hd__o21ai_2 _36003_ (.A1(_13431_),
    .A2(_13426_),
    .B1(_13428_),
    .Y(_13437_));
 sky130_fd_sc_hd__nand3_4 _36004_ (.A(_13435_),
    .B(_13436_),
    .C(_13437_),
    .Y(_13438_));
 sky130_fd_sc_hd__nor2_4 _36005_ (.A(_13252_),
    .B(_13250_),
    .Y(_13439_));
 sky130_fd_sc_hd__nor2_4 _36006_ (.A(_13251_),
    .B(_13439_),
    .Y(_13440_));
 sky130_fd_sc_hd__nand3_4 _36007_ (.A(_13434_),
    .B(_13438_),
    .C(_13440_),
    .Y(_13441_));
 sky130_fd_sc_hd__o2bb2ai_2 _36008_ (.A1_N(_13438_),
    .A2_N(_13434_),
    .B1(_13251_),
    .B2(_13439_),
    .Y(_13442_));
 sky130_fd_sc_hd__o211ai_4 _36009_ (.A1(_13425_),
    .A2(_13262_),
    .B1(_13441_),
    .C1(_13442_),
    .Y(_13443_));
 sky130_fd_sc_hd__nand2_1 _36010_ (.A(_13442_),
    .B(_13441_),
    .Y(_13444_));
 sky130_fd_sc_hd__nor2_2 _36011_ (.A(_13425_),
    .B(_13262_),
    .Y(_13445_));
 sky130_fd_sc_hd__nand2_4 _36012_ (.A(_13444_),
    .B(_13445_),
    .Y(_13446_));
 sky130_fd_sc_hd__nand3_4 _36013_ (.A(_10692_),
    .B(_06208_),
    .C(_09490_),
    .Y(_13447_));
 sky130_fd_sc_hd__nor2_4 _36014_ (.A(_10780_),
    .B(_13447_),
    .Y(_13448_));
 sky130_fd_sc_hd__nand2_2 _36015_ (.A(_19899_),
    .B(_09787_),
    .Y(_13449_));
 sky130_vsdinv _36016_ (.A(_13449_),
    .Y(_13450_));
 sky130_fd_sc_hd__buf_2 _36017_ (.A(_12102_),
    .X(_13451_));
 sky130_fd_sc_hd__a22o_2 _36018_ (.A1(_19894_),
    .A2(_13451_),
    .B1(_19897_),
    .B2(_11927_),
    .X(_13452_));
 sky130_fd_sc_hd__nand3b_4 _36019_ (.A_N(_13448_),
    .B(_13450_),
    .C(_13452_),
    .Y(_13453_));
 sky130_fd_sc_hd__a22oi_4 _36020_ (.A1(net444),
    .A2(_12109_),
    .B1(_10351_),
    .B2(_20091_),
    .Y(_13454_));
 sky130_fd_sc_hd__o21ai_4 _36021_ (.A1(_13454_),
    .A2(_13448_),
    .B1(_13449_),
    .Y(_13455_));
 sky130_fd_sc_hd__buf_4 _36022_ (.A(_09487_),
    .X(_13456_));
 sky130_fd_sc_hd__a31o_1 _36023_ (.A1(_13275_),
    .A2(net455),
    .A3(_13456_),
    .B1(_13269_),
    .X(_13457_));
 sky130_fd_sc_hd__a21oi_4 _36024_ (.A1(_13453_),
    .A2(_13455_),
    .B1(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__a21oi_4 _36025_ (.A1(_13272_),
    .A2(_13275_),
    .B1(_13269_),
    .Y(_13459_));
 sky130_fd_sc_hd__nand2_2 _36026_ (.A(_13453_),
    .B(_13455_),
    .Y(_13460_));
 sky130_fd_sc_hd__nor2_4 _36027_ (.A(_13459_),
    .B(_13460_),
    .Y(_13461_));
 sky130_fd_sc_hd__a22oi_4 _36028_ (.A1(_19903_),
    .A2(_11165_),
    .B1(_19907_),
    .B2(_20079_),
    .Y(_13462_));
 sky130_fd_sc_hd__nand2_2 _36029_ (.A(_06048_),
    .B(_20082_),
    .Y(_13463_));
 sky130_fd_sc_hd__nand2_2 _36030_ (.A(_06049_),
    .B(_20078_),
    .Y(_13464_));
 sky130_fd_sc_hd__nor2_4 _36031_ (.A(_13463_),
    .B(_13464_),
    .Y(_13465_));
 sky130_fd_sc_hd__nor2_1 _36032_ (.A(_13462_),
    .B(_13465_),
    .Y(_13466_));
 sky130_fd_sc_hd__nand2_1 _36033_ (.A(_06052_),
    .B(_20073_),
    .Y(_13467_));
 sky130_vsdinv _36034_ (.A(_13467_),
    .Y(_13468_));
 sky130_fd_sc_hd__nand2_1 _36035_ (.A(_13466_),
    .B(_13468_),
    .Y(_13469_));
 sky130_fd_sc_hd__o21ai_1 _36036_ (.A1(_13462_),
    .A2(_13465_),
    .B1(_13467_),
    .Y(_13470_));
 sky130_fd_sc_hd__nand2_2 _36037_ (.A(_13469_),
    .B(_13470_),
    .Y(_13471_));
 sky130_fd_sc_hd__o21a_1 _36038_ (.A1(_13458_),
    .A2(_13461_),
    .B1(_13471_),
    .X(_13472_));
 sky130_fd_sc_hd__o31a_1 _36039_ (.A1(_13449_),
    .A2(_13454_),
    .A3(_13448_),
    .B1(_13457_),
    .X(_13473_));
 sky130_fd_sc_hd__nand2_1 _36040_ (.A(_13473_),
    .B(_13455_),
    .Y(_13474_));
 sky130_fd_sc_hd__nand2_2 _36041_ (.A(_13460_),
    .B(_13459_),
    .Y(_13475_));
 sky130_fd_sc_hd__nand2_1 _36042_ (.A(_13466_),
    .B(_13467_),
    .Y(_13476_));
 sky130_fd_sc_hd__o21ai_1 _36043_ (.A1(_13462_),
    .A2(_13465_),
    .B1(_13468_),
    .Y(_13477_));
 sky130_fd_sc_hd__nand2_2 _36044_ (.A(_13476_),
    .B(_13477_),
    .Y(_13478_));
 sky130_fd_sc_hd__and3_1 _36045_ (.A(_13474_),
    .B(_13475_),
    .C(_13478_),
    .X(_13479_));
 sky130_fd_sc_hd__o2bb2ai_4 _36046_ (.A1_N(_13443_),
    .A2_N(_13446_),
    .B1(_13472_),
    .B2(_13479_),
    .Y(_13480_));
 sky130_fd_sc_hd__o21ai_1 _36047_ (.A1(_13458_),
    .A2(_13461_),
    .B1(_13478_),
    .Y(_13481_));
 sky130_fd_sc_hd__nand3_1 _36048_ (.A(_13474_),
    .B(_13475_),
    .C(_13471_),
    .Y(_13482_));
 sky130_fd_sc_hd__nand2_2 _36049_ (.A(_13481_),
    .B(_13482_),
    .Y(_13483_));
 sky130_fd_sc_hd__nand3_4 _36050_ (.A(_13446_),
    .B(_13483_),
    .C(_13443_),
    .Y(_13484_));
 sky130_fd_sc_hd__o21ai_4 _36051_ (.A1(_13229_),
    .A2(_13230_),
    .B1(_13223_),
    .Y(_13485_));
 sky130_fd_sc_hd__a21o_1 _36052_ (.A1(_13480_),
    .A2(_13484_),
    .B1(_13485_),
    .X(_13486_));
 sky130_fd_sc_hd__nand3_4 _36053_ (.A(_13485_),
    .B(_13480_),
    .C(_13484_),
    .Y(_13487_));
 sky130_fd_sc_hd__buf_2 _36054_ (.A(_13487_),
    .X(_13488_));
 sky130_fd_sc_hd__o21a_2 _36055_ (.A1(_13296_),
    .A2(_13264_),
    .B1(_13297_),
    .X(_13489_));
 sky130_vsdinv _36056_ (.A(_13489_),
    .Y(_13490_));
 sky130_fd_sc_hd__and3_1 _36057_ (.A(_13486_),
    .B(_13488_),
    .C(_13490_),
    .X(_13491_));
 sky130_fd_sc_hd__a21oi_4 _36058_ (.A1(_13486_),
    .A2(_13487_),
    .B1(_13490_),
    .Y(_13492_));
 sky130_fd_sc_hd__nand3_4 _36059_ (.A(_08589_),
    .B(_08591_),
    .C(_07257_),
    .Y(_13493_));
 sky130_fd_sc_hd__nor2_8 _36060_ (.A(_08040_),
    .B(_13493_),
    .Y(_13494_));
 sky130_fd_sc_hd__nand2_4 _36061_ (.A(_07967_),
    .B(_07250_),
    .Y(_13495_));
 sky130_vsdinv _36062_ (.A(_13495_),
    .Y(_13496_));
 sky130_fd_sc_hd__buf_4 _36063_ (.A(_08591_),
    .X(_13497_));
 sky130_fd_sc_hd__a22o_2 _36064_ (.A1(_12848_),
    .A2(_07543_),
    .B1(_13497_),
    .B2(_20123_),
    .X(_13498_));
 sky130_fd_sc_hd__nand3b_2 _36065_ (.A_N(_13494_),
    .B(_13496_),
    .C(_13498_),
    .Y(_13499_));
 sky130_fd_sc_hd__a21o_1 _36066_ (.A1(_13199_),
    .A2(_13197_),
    .B1(_13196_),
    .X(_13500_));
 sky130_fd_sc_hd__a22oi_4 _36067_ (.A1(_12848_),
    .A2(_07258_),
    .B1(_13497_),
    .B2(_09443_),
    .Y(_13501_));
 sky130_fd_sc_hd__o21ai_2 _36068_ (.A1(_13501_),
    .A2(_13494_),
    .B1(_13495_),
    .Y(_13502_));
 sky130_fd_sc_hd__nand3_4 _36069_ (.A(_13499_),
    .B(_13500_),
    .C(_13502_),
    .Y(_13503_));
 sky130_fd_sc_hd__o21ai_2 _36070_ (.A1(_13501_),
    .A2(_13494_),
    .B1(_13496_),
    .Y(_13504_));
 sky130_fd_sc_hd__a21oi_2 _36071_ (.A1(_13199_),
    .A2(_13197_),
    .B1(_13196_),
    .Y(_13505_));
 sky130_fd_sc_hd__o211ai_4 _36072_ (.A1(_11457_),
    .A2(_13493_),
    .B1(_13495_),
    .C1(_13498_),
    .Y(_13506_));
 sky130_fd_sc_hd__nand3_4 _36073_ (.A(_13504_),
    .B(_13505_),
    .C(_13506_),
    .Y(_13507_));
 sky130_fd_sc_hd__nand2_1 _36074_ (.A(_13503_),
    .B(_13507_),
    .Y(_13508_));
 sky130_fd_sc_hd__nand2_2 _36075_ (.A(_10934_),
    .B(_20114_),
    .Y(_13509_));
 sky130_fd_sc_hd__nand2_4 _36076_ (.A(_08248_),
    .B(_08053_),
    .Y(_13510_));
 sky130_fd_sc_hd__nor2_4 _36077_ (.A(_13509_),
    .B(_13510_),
    .Y(_13511_));
 sky130_fd_sc_hd__and2_1 _36078_ (.A(_13509_),
    .B(_13510_),
    .X(_13512_));
 sky130_fd_sc_hd__nand2_1 _36079_ (.A(_11869_),
    .B(_11723_),
    .Y(_13513_));
 sky130_fd_sc_hd__o21bai_4 _36080_ (.A1(_13511_),
    .A2(_13512_),
    .B1_N(_13513_),
    .Y(_13514_));
 sky130_fd_sc_hd__nand3_1 _36081_ (.A(_07483_),
    .B(_11871_),
    .C(_10711_),
    .Y(_13515_));
 sky130_fd_sc_hd__nand2_1 _36082_ (.A(_13509_),
    .B(_13510_),
    .Y(_13516_));
 sky130_fd_sc_hd__o211a_1 _36083_ (.A1(_11057_),
    .A2(_13515_),
    .B1(_13513_),
    .C1(_13516_),
    .X(_13517_));
 sky130_vsdinv _36084_ (.A(_13517_),
    .Y(_13518_));
 sky130_fd_sc_hd__nand3_4 _36085_ (.A(_13508_),
    .B(_13514_),
    .C(_13518_),
    .Y(_13519_));
 sky130_fd_sc_hd__nand2_2 _36086_ (.A(_13518_),
    .B(_13514_),
    .Y(_13520_));
 sky130_fd_sc_hd__nand3_4 _36087_ (.A(_13520_),
    .B(_13503_),
    .C(_13507_),
    .Y(_13521_));
 sky130_fd_sc_hd__nand2_1 _36088_ (.A(_13133_),
    .B(_13130_),
    .Y(_13522_));
 sky130_fd_sc_hd__nand2_4 _36089_ (.A(_13522_),
    .B(_13126_),
    .Y(_13523_));
 sky130_fd_sc_hd__a21o_2 _36090_ (.A1(_13519_),
    .A2(_13521_),
    .B1(_13523_),
    .X(_13524_));
 sky130_fd_sc_hd__nand3_1 _36091_ (.A(_13523_),
    .B(_13519_),
    .C(_13521_),
    .Y(_13525_));
 sky130_fd_sc_hd__buf_2 _36092_ (.A(_13525_),
    .X(_13526_));
 sky130_fd_sc_hd__nand2_1 _36093_ (.A(_13214_),
    .B(_13206_),
    .Y(_13527_));
 sky130_fd_sc_hd__nand2_4 _36094_ (.A(_13527_),
    .B(_13203_),
    .Y(_13528_));
 sky130_fd_sc_hd__a21oi_4 _36095_ (.A1(_13524_),
    .A2(_13526_),
    .B1(_13528_),
    .Y(_13529_));
 sky130_fd_sc_hd__and3_1 _36096_ (.A(_13524_),
    .B(_13526_),
    .C(_13528_),
    .X(_13530_));
 sky130_fd_sc_hd__nand2_2 _36097_ (.A(_10552_),
    .B(_06312_),
    .Y(_13531_));
 sky130_fd_sc_hd__nand2_2 _36098_ (.A(_10553_),
    .B(_08546_),
    .Y(_13532_));
 sky130_fd_sc_hd__nor2_4 _36099_ (.A(_13531_),
    .B(_13532_),
    .Y(_13533_));
 sky130_fd_sc_hd__and2_1 _36100_ (.A(_13531_),
    .B(_13532_),
    .X(_13534_));
 sky130_fd_sc_hd__nand2_2 _36101_ (.A(_19854_),
    .B(_12846_),
    .Y(_13535_));
 sky130_fd_sc_hd__o21ai_2 _36102_ (.A1(_13533_),
    .A2(_13534_),
    .B1(_13535_),
    .Y(_13536_));
 sky130_fd_sc_hd__or2_1 _36103_ (.A(_13531_),
    .B(_13532_),
    .X(_13537_));
 sky130_fd_sc_hd__nand2_2 _36104_ (.A(_13531_),
    .B(_13532_),
    .Y(_13538_));
 sky130_vsdinv _36105_ (.A(_13535_),
    .Y(_13539_));
 sky130_fd_sc_hd__nand3_2 _36106_ (.A(_13537_),
    .B(_13538_),
    .C(_13539_),
    .Y(_13540_));
 sky130_fd_sc_hd__a21o_1 _36107_ (.A1(_13163_),
    .A2(_13164_),
    .B1(_13162_),
    .X(_13541_));
 sky130_fd_sc_hd__nand3_4 _36108_ (.A(_13536_),
    .B(_13540_),
    .C(_13541_),
    .Y(_13542_));
 sky130_fd_sc_hd__o21ai_2 _36109_ (.A1(_13533_),
    .A2(_13534_),
    .B1(_13539_),
    .Y(_13543_));
 sky130_fd_sc_hd__nand3_2 _36110_ (.A(_13537_),
    .B(_13538_),
    .C(_13535_),
    .Y(_13544_));
 sky130_fd_sc_hd__a21oi_4 _36111_ (.A1(_13163_),
    .A2(_13164_),
    .B1(_13162_),
    .Y(_13545_));
 sky130_fd_sc_hd__nand3_4 _36112_ (.A(_13543_),
    .B(_13544_),
    .C(_13545_),
    .Y(_13546_));
 sky130_fd_sc_hd__a21oi_4 _36113_ (.A1(_13122_),
    .A2(_13120_),
    .B1(_13119_),
    .Y(_13547_));
 sky130_vsdinv _36114_ (.A(_13547_),
    .Y(_13548_));
 sky130_fd_sc_hd__a21oi_4 _36115_ (.A1(_13542_),
    .A2(_13546_),
    .B1(_13548_),
    .Y(_13549_));
 sky130_fd_sc_hd__nand2_2 _36116_ (.A(_13542_),
    .B(_13546_),
    .Y(_13550_));
 sky130_fd_sc_hd__nor2_4 _36117_ (.A(_13547_),
    .B(_13550_),
    .Y(_13551_));
 sky130_fd_sc_hd__nand2_2 _36118_ (.A(_11794_),
    .B(_05835_),
    .Y(_13552_));
 sky130_fd_sc_hd__nand2_2 _36119_ (.A(_10989_),
    .B(_05999_),
    .Y(_13553_));
 sky130_fd_sc_hd__nor2_4 _36120_ (.A(_13552_),
    .B(_13553_),
    .Y(_13554_));
 sky130_fd_sc_hd__nand2_2 _36121_ (.A(_19843_),
    .B(_07502_),
    .Y(_13555_));
 sky130_vsdinv _36122_ (.A(_13555_),
    .Y(_13556_));
 sky130_fd_sc_hd__nand2_1 _36123_ (.A(_13552_),
    .B(_13553_),
    .Y(_13557_));
 sky130_fd_sc_hd__nand2_2 _36124_ (.A(_13556_),
    .B(_13557_),
    .Y(_13558_));
 sky130_fd_sc_hd__nor2_2 _36125_ (.A(_13554_),
    .B(_13558_),
    .Y(_13559_));
 sky130_fd_sc_hd__and2_1 _36126_ (.A(_13552_),
    .B(_13553_),
    .X(_13560_));
 sky130_fd_sc_hd__o21ai_1 _36127_ (.A1(_13554_),
    .A2(_13560_),
    .B1(_13555_),
    .Y(_13561_));
 sky130_vsdinv _36128_ (.A(_13561_),
    .Y(_13562_));
 sky130_fd_sc_hd__o21ai_2 _36129_ (.A1(_13141_),
    .A2(_13147_),
    .B1(_13144_),
    .Y(_13563_));
 sky130_fd_sc_hd__nand3_2 _36130_ (.A(_18694_),
    .B(_13138_),
    .C(_05832_),
    .Y(_13564_));
 sky130_fd_sc_hd__nor2_2 _36131_ (.A(_20157_),
    .B(_13564_),
    .Y(_13565_));
 sky130_fd_sc_hd__a22oi_4 _36132_ (.A1(_12492_),
    .A2(_05979_),
    .B1(net446),
    .B2(_13139_),
    .Y(_13566_));
 sky130_fd_sc_hd__o22ai_4 _36133_ (.A1(_10404_),
    .A2(_06004_),
    .B1(_13565_),
    .B2(_13566_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand2_1 _36134_ (.A(_11783_),
    .B(_20152_),
    .Y(_13568_));
 sky130_fd_sc_hd__nand3b_4 _36135_ (.A_N(_13568_),
    .B(_18694_),
    .C(_06256_),
    .Y(_13569_));
 sky130_fd_sc_hd__o21ai_2 _36136_ (.A1(_20157_),
    .A2(_11275_),
    .B1(_13568_),
    .Y(_13570_));
 sky130_fd_sc_hd__nand2_2 _36137_ (.A(_19833_),
    .B(_06148_),
    .Y(_13571_));
 sky130_vsdinv _36138_ (.A(_13571_),
    .Y(_13572_));
 sky130_fd_sc_hd__nand3_4 _36139_ (.A(_13569_),
    .B(_13570_),
    .C(_13572_),
    .Y(_13573_));
 sky130_fd_sc_hd__a22oi_4 _36140_ (.A1(_13148_),
    .A2(_13563_),
    .B1(_13567_),
    .B2(_13573_),
    .Y(_13574_));
 sky130_fd_sc_hd__a21oi_4 _36141_ (.A1(_13147_),
    .A2(_13141_),
    .B1(_13144_),
    .Y(_13575_));
 sky130_fd_sc_hd__o211a_1 _36142_ (.A1(_13143_),
    .A2(_13575_),
    .B1(_13573_),
    .C1(_13567_),
    .X(_13576_));
 sky130_fd_sc_hd__o22ai_4 _36143_ (.A1(_13559_),
    .A2(_13562_),
    .B1(_13574_),
    .B2(_13576_),
    .Y(_13577_));
 sky130_fd_sc_hd__o21a_1 _36144_ (.A1(_13141_),
    .A2(_13147_),
    .B1(_13144_),
    .X(_13578_));
 sky130_fd_sc_hd__o21bai_1 _36145_ (.A1(_20157_),
    .A2(_13564_),
    .B1_N(_13571_),
    .Y(_13579_));
 sky130_fd_sc_hd__nor2_2 _36146_ (.A(_13566_),
    .B(_13579_),
    .Y(_13580_));
 sky130_fd_sc_hd__a21oi_2 _36147_ (.A1(_13569_),
    .A2(_13570_),
    .B1(_13572_),
    .Y(_13581_));
 sky130_fd_sc_hd__o22ai_4 _36148_ (.A1(_13140_),
    .A2(_13578_),
    .B1(_13580_),
    .B2(_13581_),
    .Y(_13582_));
 sky130_fd_sc_hd__o211ai_4 _36149_ (.A1(_13143_),
    .A2(_13575_),
    .B1(_13573_),
    .C1(_13567_),
    .Y(_13583_));
 sky130_fd_sc_hd__o21ai_1 _36150_ (.A1(_13554_),
    .A2(_13560_),
    .B1(_13556_),
    .Y(_13584_));
 sky130_fd_sc_hd__or2_2 _36151_ (.A(_13552_),
    .B(_13553_),
    .X(_13585_));
 sky130_fd_sc_hd__nand3_1 _36152_ (.A(_13585_),
    .B(_13557_),
    .C(_13555_),
    .Y(_13586_));
 sky130_fd_sc_hd__nand2_2 _36153_ (.A(_13584_),
    .B(_13586_),
    .Y(_13587_));
 sky130_fd_sc_hd__nand3_4 _36154_ (.A(_13582_),
    .B(_13583_),
    .C(_13587_),
    .Y(_13588_));
 sky130_fd_sc_hd__nand2_1 _36155_ (.A(_13152_),
    .B(_13171_),
    .Y(_13589_));
 sky130_fd_sc_hd__nand2_4 _36156_ (.A(_13589_),
    .B(_13156_),
    .Y(_13590_));
 sky130_fd_sc_hd__a21oi_4 _36157_ (.A1(_13577_),
    .A2(_13588_),
    .B1(_13590_),
    .Y(_13591_));
 sky130_fd_sc_hd__and3_1 _36158_ (.A(_13153_),
    .B(_13154_),
    .C(_13155_),
    .X(_13592_));
 sky130_fd_sc_hd__a31oi_1 _36159_ (.A1(_13146_),
    .A2(_13150_),
    .A3(_13151_),
    .B1(_13179_),
    .Y(_13593_));
 sky130_fd_sc_hd__o211a_2 _36160_ (.A1(_13592_),
    .A2(_13593_),
    .B1(_13588_),
    .C1(_13577_),
    .X(_13594_));
 sky130_fd_sc_hd__o22ai_4 _36161_ (.A1(_13549_),
    .A2(_13551_),
    .B1(_13591_),
    .B2(_13594_),
    .Y(_13595_));
 sky130_fd_sc_hd__a21o_1 _36162_ (.A1(_13577_),
    .A2(_13588_),
    .B1(_13590_),
    .X(_13596_));
 sky130_fd_sc_hd__nor2_4 _36163_ (.A(_13549_),
    .B(_13551_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand3_4 _36164_ (.A(_13590_),
    .B(_13577_),
    .C(_13588_),
    .Y(_13598_));
 sky130_fd_sc_hd__nand3_4 _36165_ (.A(_13596_),
    .B(_13597_),
    .C(_13598_),
    .Y(_13599_));
 sky130_fd_sc_hd__nand2_2 _36166_ (.A(_13137_),
    .B(_13181_),
    .Y(_13600_));
 sky130_fd_sc_hd__nand2_2 _36167_ (.A(_13600_),
    .B(_13173_),
    .Y(_13601_));
 sky130_fd_sc_hd__a21oi_4 _36168_ (.A1(_13595_),
    .A2(_13599_),
    .B1(_13601_),
    .Y(_13602_));
 sky130_vsdinv _36169_ (.A(_13173_),
    .Y(_13603_));
 sky130_fd_sc_hd__a31oi_4 _36170_ (.A1(_13178_),
    .A2(_13180_),
    .A3(_13177_),
    .B1(_13190_),
    .Y(_13604_));
 sky130_fd_sc_hd__o211a_1 _36171_ (.A1(_13603_),
    .A2(_13604_),
    .B1(_13599_),
    .C1(_13595_),
    .X(_13605_));
 sky130_fd_sc_hd__o22ai_4 _36172_ (.A1(_13529_),
    .A2(_13530_),
    .B1(_13602_),
    .B2(_13605_),
    .Y(_13606_));
 sky130_fd_sc_hd__nand2_1 _36173_ (.A(_13595_),
    .B(_13599_),
    .Y(_13607_));
 sky130_fd_sc_hd__nor2_1 _36174_ (.A(_13603_),
    .B(_13604_),
    .Y(_13608_));
 sky130_fd_sc_hd__nand2_1 _36175_ (.A(_13607_),
    .B(_13608_),
    .Y(_13609_));
 sky130_fd_sc_hd__nand3_4 _36176_ (.A(_13601_),
    .B(_13595_),
    .C(_13599_),
    .Y(_13610_));
 sky130_vsdinv _36177_ (.A(_13528_),
    .Y(_13611_));
 sky130_fd_sc_hd__a21o_1 _36178_ (.A1(_13524_),
    .A2(_13526_),
    .B1(_13611_),
    .X(_13612_));
 sky130_fd_sc_hd__nand3_1 _36179_ (.A(_13524_),
    .B(_13526_),
    .C(_13611_),
    .Y(_13613_));
 sky130_fd_sc_hd__nand2_1 _36180_ (.A(_13612_),
    .B(_13613_),
    .Y(_13614_));
 sky130_fd_sc_hd__nand3_4 _36181_ (.A(_13609_),
    .B(_13610_),
    .C(_13614_),
    .Y(_13615_));
 sky130_fd_sc_hd__nand2_2 _36182_ (.A(_13183_),
    .B(_13182_),
    .Y(_13616_));
 sky130_fd_sc_hd__nor2_4 _36183_ (.A(_13187_),
    .B(_13616_),
    .Y(_13617_));
 sky130_fd_sc_hd__a21o_2 _36184_ (.A1(_13232_),
    .A2(_13192_),
    .B1(_13617_),
    .X(_13618_));
 sky130_fd_sc_hd__a21oi_4 _36185_ (.A1(_13606_),
    .A2(_13615_),
    .B1(_13618_),
    .Y(_13619_));
 sky130_fd_sc_hd__a21oi_4 _36186_ (.A1(_13187_),
    .A2(_13616_),
    .B1(_13239_),
    .Y(_13620_));
 sky130_fd_sc_hd__o211a_2 _36187_ (.A1(_13617_),
    .A2(_13620_),
    .B1(_13615_),
    .C1(_13606_),
    .X(_13621_));
 sky130_fd_sc_hd__o22ai_4 _36188_ (.A1(_13491_),
    .A2(_13492_),
    .B1(_13619_),
    .B2(_13621_),
    .Y(_13622_));
 sky130_fd_sc_hd__a21bo_1 _36189_ (.A1(_13312_),
    .A2(_13241_),
    .B1_N(_13234_),
    .X(_13623_));
 sky130_fd_sc_hd__a21o_1 _36190_ (.A1(_13606_),
    .A2(_13615_),
    .B1(_13618_),
    .X(_13624_));
 sky130_fd_sc_hd__a21oi_4 _36191_ (.A1(_13480_),
    .A2(_13484_),
    .B1(_13485_),
    .Y(_13625_));
 sky130_fd_sc_hd__nor2_2 _36192_ (.A(_13489_),
    .B(_13625_),
    .Y(_13626_));
 sky130_fd_sc_hd__a21oi_4 _36193_ (.A1(_13488_),
    .A2(_13626_),
    .B1(_13492_),
    .Y(_13627_));
 sky130_fd_sc_hd__nand3_4 _36194_ (.A(_13618_),
    .B(_13606_),
    .C(_13615_),
    .Y(_13628_));
 sky130_fd_sc_hd__nand3_2 _36195_ (.A(_13624_),
    .B(_13627_),
    .C(_13628_),
    .Y(_13629_));
 sky130_fd_sc_hd__nand3_4 _36196_ (.A(_13622_),
    .B(_13623_),
    .C(_13629_),
    .Y(_13630_));
 sky130_fd_sc_hd__o21ai_2 _36197_ (.A1(_13619_),
    .A2(_13621_),
    .B1(_13627_),
    .Y(_13631_));
 sky130_fd_sc_hd__a21boi_2 _36198_ (.A1(_13312_),
    .A2(_13241_),
    .B1_N(_13234_),
    .Y(_13632_));
 sky130_fd_sc_hd__a21o_1 _36199_ (.A1(_13486_),
    .A2(_13488_),
    .B1(_13490_),
    .X(_13633_));
 sky130_fd_sc_hd__nand2_1 _36200_ (.A(_13626_),
    .B(_13488_),
    .Y(_13634_));
 sky130_fd_sc_hd__nand2_2 _36201_ (.A(_13633_),
    .B(_13634_),
    .Y(_13635_));
 sky130_fd_sc_hd__nand3_2 _36202_ (.A(_13624_),
    .B(_13628_),
    .C(_13635_),
    .Y(_13636_));
 sky130_fd_sc_hd__nand3_4 _36203_ (.A(_13631_),
    .B(_13632_),
    .C(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__nand2_2 _36204_ (.A(_10809_),
    .B(_20069_),
    .Y(_13638_));
 sky130_fd_sc_hd__nand2_2 _36205_ (.A(_18686_),
    .B(_06098_),
    .Y(_13639_));
 sky130_fd_sc_hd__nor2_4 _36206_ (.A(_13638_),
    .B(_13639_),
    .Y(_13640_));
 sky130_fd_sc_hd__and2_1 _36207_ (.A(_13638_),
    .B(_13639_),
    .X(_13641_));
 sky130_fd_sc_hd__o21ai_2 _36208_ (.A1(_13640_),
    .A2(_13641_),
    .B1(_13329_),
    .Y(_13642_));
 sky130_fd_sc_hd__or2_1 _36209_ (.A(_13638_),
    .B(_13639_),
    .X(_13643_));
 sky130_fd_sc_hd__nand2_2 _36210_ (.A(_13638_),
    .B(_13639_),
    .Y(_13644_));
 sky130_fd_sc_hd__nand3_2 _36211_ (.A(_13643_),
    .B(_13325_),
    .C(_13644_),
    .Y(_13645_));
 sky130_fd_sc_hd__nand2_2 _36212_ (.A(_13281_),
    .B(_13282_),
    .Y(_13646_));
 sky130_fd_sc_hd__buf_6 _36213_ (.A(_10761_),
    .X(_13647_));
 sky130_fd_sc_hd__a31o_1 _36214_ (.A1(_13646_),
    .A2(_19910_),
    .A3(_13647_),
    .B1(_13283_),
    .X(_13648_));
 sky130_fd_sc_hd__nand3_4 _36215_ (.A(_13642_),
    .B(_13645_),
    .C(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__o21ai_2 _36216_ (.A1(_13640_),
    .A2(_13641_),
    .B1(_13325_),
    .Y(_13650_));
 sky130_fd_sc_hd__nand3_2 _36217_ (.A(_13643_),
    .B(_13329_),
    .C(_13644_),
    .Y(_13651_));
 sky130_fd_sc_hd__a21oi_4 _36218_ (.A1(_13285_),
    .A2(_13646_),
    .B1(_13283_),
    .Y(_13652_));
 sky130_fd_sc_hd__nand3_4 _36219_ (.A(_13650_),
    .B(_13651_),
    .C(_13652_),
    .Y(_13653_));
 sky130_fd_sc_hd__nor2_4 _36220_ (.A(_13325_),
    .B(_13322_),
    .Y(_13654_));
 sky130_fd_sc_hd__o2bb2ai_4 _36221_ (.A1_N(_13649_),
    .A2_N(_13653_),
    .B1(_13320_),
    .B2(_13654_),
    .Y(_13655_));
 sky130_fd_sc_hd__nor2_4 _36222_ (.A(_13320_),
    .B(_13654_),
    .Y(_13656_));
 sky130_fd_sc_hd__nand3_4 _36223_ (.A(_13649_),
    .B(_13653_),
    .C(_13656_),
    .Y(_13657_));
 sky130_fd_sc_hd__nand2_1 _36224_ (.A(_13655_),
    .B(_13657_),
    .Y(_13658_));
 sky130_fd_sc_hd__o21a_1 _36225_ (.A1(_13288_),
    .A2(_13290_),
    .B1(_13277_),
    .X(_13659_));
 sky130_fd_sc_hd__nand2_2 _36226_ (.A(_13658_),
    .B(_13659_),
    .Y(_13660_));
 sky130_fd_sc_hd__o21ai_4 _36227_ (.A1(_13288_),
    .A2(_13290_),
    .B1(_13277_),
    .Y(_13661_));
 sky130_fd_sc_hd__nand3_4 _36228_ (.A(_13661_),
    .B(_13655_),
    .C(_13657_),
    .Y(_13662_));
 sky130_fd_sc_hd__and2_2 _36229_ (.A(_13345_),
    .B(_13336_),
    .X(_13663_));
 sky130_fd_sc_hd__a21o_1 _36230_ (.A1(_13660_),
    .A2(_13662_),
    .B1(_13663_),
    .X(_13664_));
 sky130_fd_sc_hd__nand2_1 _36231_ (.A(_13353_),
    .B(_13352_),
    .Y(_13665_));
 sky130_fd_sc_hd__nand2_1 _36232_ (.A(_13665_),
    .B(_13351_),
    .Y(_13666_));
 sky130_fd_sc_hd__nand3_2 _36233_ (.A(_13660_),
    .B(_13663_),
    .C(_13662_),
    .Y(_13667_));
 sky130_fd_sc_hd__nand3_4 _36234_ (.A(_13664_),
    .B(_13666_),
    .C(_13667_),
    .Y(_13668_));
 sky130_fd_sc_hd__a21bo_1 _36235_ (.A1(_13660_),
    .A2(_13662_),
    .B1_N(_13663_),
    .X(_13669_));
 sky130_fd_sc_hd__and2_1 _36236_ (.A(_13665_),
    .B(_13351_),
    .X(_13670_));
 sky130_fd_sc_hd__nand3b_2 _36237_ (.A_N(_13663_),
    .B(_13660_),
    .C(_13662_),
    .Y(_13671_));
 sky130_fd_sc_hd__nand3_4 _36238_ (.A(_13669_),
    .B(_13670_),
    .C(_13671_),
    .Y(_13672_));
 sky130_fd_sc_hd__and3_1 _36239_ (.A(_11603_),
    .B(_19921_),
    .C(_19926_),
    .X(_13673_));
 sky130_fd_sc_hd__nand3_4 _36240_ (.A(_12355_),
    .B(_19939_),
    .C(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__a21oi_4 _36241_ (.A1(_13367_),
    .A2(_13674_),
    .B1(_12673_),
    .Y(_13675_));
 sky130_fd_sc_hd__and3_2 _36242_ (.A(_13367_),
    .B(_12673_),
    .C(_13674_),
    .X(_13676_));
 sky130_fd_sc_hd__nor2_8 _36243_ (.A(_13675_),
    .B(_13676_),
    .Y(_13677_));
 sky130_vsdinv _36244_ (.A(_13677_),
    .Y(_13678_));
 sky130_fd_sc_hd__buf_4 _36245_ (.A(_13678_),
    .X(_13679_));
 sky130_fd_sc_hd__a21o_1 _36246_ (.A1(_13668_),
    .A2(_13672_),
    .B1(_13679_),
    .X(_13680_));
 sky130_fd_sc_hd__a21oi_4 _36247_ (.A1(_13293_),
    .A2(_13298_),
    .B1(_13294_),
    .Y(_13681_));
 sky130_fd_sc_hd__a21oi_4 _36248_ (.A1(_13299_),
    .A2(_13305_),
    .B1(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__nand3_4 _36249_ (.A(_13672_),
    .B(_13668_),
    .C(_13679_),
    .Y(_13683_));
 sky130_fd_sc_hd__nand3_4 _36250_ (.A(_13680_),
    .B(_13682_),
    .C(_13683_),
    .Y(_13684_));
 sky130_fd_sc_hd__a31oi_4 _36251_ (.A1(_13293_),
    .A2(_13298_),
    .A3(_13294_),
    .B1(_13310_),
    .Y(_13685_));
 sky130_fd_sc_hd__buf_2 _36252_ (.A(_13677_),
    .X(_13686_));
 sky130_fd_sc_hd__buf_4 _36253_ (.A(_13686_),
    .X(_13687_));
 sky130_fd_sc_hd__nand3_2 _36254_ (.A(_13672_),
    .B(_13668_),
    .C(_13687_),
    .Y(_13688_));
 sky130_fd_sc_hd__buf_6 _36255_ (.A(_13676_),
    .X(_13689_));
 sky130_fd_sc_hd__o2bb2ai_2 _36256_ (.A1_N(_13668_),
    .A2_N(_13672_),
    .B1(_13689_),
    .B2(_13675_),
    .Y(_13690_));
 sky130_fd_sc_hd__o211ai_4 _36257_ (.A1(_13681_),
    .A2(_13685_),
    .B1(_13688_),
    .C1(_13690_),
    .Y(_13691_));
 sky130_vsdinv _36258_ (.A(_13361_),
    .Y(_13692_));
 sky130_fd_sc_hd__and2_1 _36259_ (.A(_13355_),
    .B(_13369_),
    .X(_13693_));
 sky130_fd_sc_hd__nor2_4 _36260_ (.A(_13692_),
    .B(_13693_),
    .Y(_13694_));
 sky130_vsdinv _36261_ (.A(_13694_),
    .Y(_13695_));
 sky130_fd_sc_hd__a21oi_4 _36262_ (.A1(_13684_),
    .A2(_13691_),
    .B1(_13695_),
    .Y(_13696_));
 sky130_fd_sc_hd__and3_1 _36263_ (.A(_13695_),
    .B(_13684_),
    .C(_13691_),
    .X(_13697_));
 sky130_fd_sc_hd__o2bb2ai_2 _36264_ (.A1_N(_13630_),
    .A2_N(_13637_),
    .B1(_13696_),
    .B2(_13697_),
    .Y(_13698_));
 sky130_fd_sc_hd__a21bo_1 _36265_ (.A1(_13386_),
    .A2(_13319_),
    .B1_N(_13314_),
    .X(_13699_));
 sky130_fd_sc_hd__a31oi_4 _36266_ (.A1(_13680_),
    .A2(_13682_),
    .A3(_13683_),
    .B1(_13694_),
    .Y(_13700_));
 sky130_fd_sc_hd__a21oi_4 _36267_ (.A1(_13691_),
    .A2(_13700_),
    .B1(_13696_),
    .Y(_13701_));
 sky130_fd_sc_hd__nand3_2 _36268_ (.A(_13637_),
    .B(_13701_),
    .C(_13630_),
    .Y(_13702_));
 sky130_fd_sc_hd__nand3_4 _36269_ (.A(_13698_),
    .B(_13699_),
    .C(_13702_),
    .Y(_13703_));
 sky130_fd_sc_hd__nand2_1 _36270_ (.A(_13637_),
    .B(_13630_),
    .Y(_13704_));
 sky130_fd_sc_hd__nand2_1 _36271_ (.A(_13704_),
    .B(_13701_),
    .Y(_13705_));
 sky130_fd_sc_hd__a21boi_2 _36272_ (.A1(_13386_),
    .A2(_13319_),
    .B1_N(_13314_),
    .Y(_13706_));
 sky130_fd_sc_hd__o211ai_4 _36273_ (.A1(_13696_),
    .A2(_13697_),
    .B1(_13630_),
    .C1(_13637_),
    .Y(_13707_));
 sky130_fd_sc_hd__nand3_4 _36274_ (.A(_13705_),
    .B(_13706_),
    .C(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__nand2_1 _36275_ (.A(_13368_),
    .B(_13674_),
    .Y(_13709_));
 sky130_fd_sc_hd__and2_2 _36276_ (.A(_13382_),
    .B(_13375_),
    .X(_13710_));
 sky130_fd_sc_hd__nor2_1 _36277_ (.A(_13709_),
    .B(_13710_),
    .Y(_13711_));
 sky130_fd_sc_hd__and3_1 _36278_ (.A(_13382_),
    .B(_13375_),
    .C(_13709_),
    .X(_13712_));
 sky130_fd_sc_hd__o2bb2ai_2 _36279_ (.A1_N(_13703_),
    .A2_N(_13708_),
    .B1(_13711_),
    .B2(_13712_),
    .Y(_13713_));
 sky130_fd_sc_hd__o21a_1 _36280_ (.A1(_13401_),
    .A2(_13389_),
    .B1(_13400_),
    .X(_13714_));
 sky130_vsdinv _36281_ (.A(_13709_),
    .Y(_13715_));
 sky130_fd_sc_hd__and3_1 _36282_ (.A(_13382_),
    .B(_13375_),
    .C(_13715_),
    .X(_13716_));
 sky130_fd_sc_hd__nor2_8 _36283_ (.A(_13715_),
    .B(_13710_),
    .Y(_13717_));
 sky130_fd_sc_hd__nor2_4 _36284_ (.A(_13716_),
    .B(_13717_),
    .Y(_13718_));
 sky130_fd_sc_hd__nand3b_2 _36285_ (.A_N(_13718_),
    .B(_13708_),
    .C(_13703_),
    .Y(_13719_));
 sky130_fd_sc_hd__nand3_4 _36286_ (.A(_13713_),
    .B(_13714_),
    .C(_13719_),
    .Y(_13720_));
 sky130_fd_sc_hd__o2bb2ai_2 _36287_ (.A1_N(_13703_),
    .A2_N(_13708_),
    .B1(_13717_),
    .B2(_13716_),
    .Y(_13721_));
 sky130_fd_sc_hd__nand3_2 _36288_ (.A(_13708_),
    .B(_13703_),
    .C(_13718_),
    .Y(_13722_));
 sky130_fd_sc_hd__o21ai_2 _36289_ (.A1(_13401_),
    .A2(_13389_),
    .B1(_13400_),
    .Y(_13723_));
 sky130_fd_sc_hd__nand3_4 _36290_ (.A(_13721_),
    .B(_13722_),
    .C(_13723_),
    .Y(_13724_));
 sky130_fd_sc_hd__a21oi_4 _36291_ (.A1(_13720_),
    .A2(_13724_),
    .B1(_13405_),
    .Y(_13725_));
 sky130_fd_sc_hd__and3_1 _36292_ (.A(_13407_),
    .B(_13409_),
    .C(_13408_),
    .X(_13726_));
 sky130_fd_sc_hd__a31oi_4 _36293_ (.A1(_13102_),
    .A2(_13398_),
    .A3(_13402_),
    .B1(_13072_),
    .Y(_13727_));
 sky130_fd_sc_hd__nand3_2 _36294_ (.A(_13720_),
    .B(_13724_),
    .C(_13405_),
    .Y(_13728_));
 sky130_fd_sc_hd__o21ai_4 _36295_ (.A1(_13726_),
    .A2(_13727_),
    .B1(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__nand2_1 _36296_ (.A(_13720_),
    .B(_13724_),
    .Y(_13730_));
 sky130_fd_sc_hd__nand2_1 _36297_ (.A(_13730_),
    .B(_13405_),
    .Y(_13731_));
 sky130_fd_sc_hd__nand3b_2 _36298_ (.A_N(_13405_),
    .B(_13720_),
    .C(_13724_),
    .Y(_13732_));
 sky130_fd_sc_hd__a21boi_2 _36299_ (.A1(_13403_),
    .A2(_13082_),
    .B1_N(_13410_),
    .Y(_13733_));
 sky130_fd_sc_hd__nand3_4 _36300_ (.A(_13731_),
    .B(_13732_),
    .C(_13733_),
    .Y(_13734_));
 sky130_fd_sc_hd__o21a_2 _36301_ (.A1(_13725_),
    .A2(_13729_),
    .B1(_13734_),
    .X(_13735_));
 sky130_fd_sc_hd__o211a_1 _36302_ (.A1(_13413_),
    .A2(_13096_),
    .B1(_13416_),
    .C1(_13417_),
    .X(_13736_));
 sky130_fd_sc_hd__a21oi_4 _36303_ (.A1(_13424_),
    .A2(_13415_),
    .B1(_13736_),
    .Y(_13737_));
 sky130_fd_sc_hd__xnor2_4 _36304_ (.A(_13735_),
    .B(_13737_),
    .Y(_02658_));
 sky130_vsdinv _36305_ (.A(_13674_),
    .Y(_13738_));
 sky130_fd_sc_hd__nor2_8 _36306_ (.A(_13738_),
    .B(_13689_),
    .Y(_13739_));
 sky130_fd_sc_hd__buf_6 _36307_ (.A(_13739_),
    .X(_13740_));
 sky130_vsdinv _36308_ (.A(_13691_),
    .Y(_13741_));
 sky130_fd_sc_hd__nor2_2 _36309_ (.A(_13700_),
    .B(_13741_),
    .Y(_13742_));
 sky130_fd_sc_hd__nor2_1 _36310_ (.A(_13740_),
    .B(_13742_),
    .Y(_13743_));
 sky130_fd_sc_hd__buf_2 _36311_ (.A(_13743_),
    .X(_13744_));
 sky130_fd_sc_hd__and2_1 _36312_ (.A(_13742_),
    .B(_13739_),
    .X(_13745_));
 sky130_fd_sc_hd__o21ai_2 _36313_ (.A1(_13635_),
    .A2(_13619_),
    .B1(_13628_),
    .Y(_13746_));
 sky130_fd_sc_hd__nand2_2 _36314_ (.A(_10067_),
    .B(_09476_),
    .Y(_13747_));
 sky130_fd_sc_hd__a21o_1 _36315_ (.A1(_19888_),
    .A2(_12304_),
    .B1(_13747_),
    .X(_13748_));
 sky130_fd_sc_hd__nand2_1 _36316_ (.A(_19887_),
    .B(_11503_),
    .Y(_13749_));
 sky130_fd_sc_hd__a21o_1 _36317_ (.A1(_19882_),
    .A2(_12303_),
    .B1(_13749_),
    .X(_13750_));
 sky130_fd_sc_hd__nand2_2 _36318_ (.A(_19890_),
    .B(_09490_),
    .Y(_13751_));
 sky130_fd_sc_hd__nand3_4 _36319_ (.A(_13748_),
    .B(_13750_),
    .C(_13751_),
    .Y(_13752_));
 sky130_fd_sc_hd__nand3b_4 _36320_ (.A_N(_13747_),
    .B(_06638_),
    .C(_09493_),
    .Y(_13753_));
 sky130_vsdinv _36321_ (.A(_13751_),
    .Y(_13754_));
 sky130_fd_sc_hd__nand2_1 _36322_ (.A(_13747_),
    .B(_13749_),
    .Y(_13755_));
 sky130_fd_sc_hd__nand3_2 _36323_ (.A(_13753_),
    .B(_13754_),
    .C(_13755_),
    .Y(_13756_));
 sky130_fd_sc_hd__clkbuf_4 _36324_ (.A(_13756_),
    .X(_13757_));
 sky130_fd_sc_hd__buf_4 _36325_ (.A(_11723_),
    .X(_13758_));
 sky130_fd_sc_hd__a31o_2 _36326_ (.A1(_13516_),
    .A2(_19879_),
    .A3(_13758_),
    .B1(_13511_),
    .X(_13759_));
 sky130_fd_sc_hd__a21oi_4 _36327_ (.A1(_13752_),
    .A2(_13757_),
    .B1(_13759_),
    .Y(_13760_));
 sky130_fd_sc_hd__a21oi_2 _36328_ (.A1(_13509_),
    .A2(_13510_),
    .B1(_13513_),
    .Y(_13761_));
 sky130_fd_sc_hd__o211a_1 _36329_ (.A1(_13511_),
    .A2(_13761_),
    .B1(_13757_),
    .C1(_13752_),
    .X(_13762_));
 sky130_fd_sc_hd__a21o_2 _36330_ (.A1(_13427_),
    .A2(_13432_),
    .B1(_13426_),
    .X(_13763_));
 sky130_fd_sc_hd__o21ai_2 _36331_ (.A1(_13760_),
    .A2(_13762_),
    .B1(_13763_),
    .Y(_13764_));
 sky130_fd_sc_hd__a21boi_2 _36332_ (.A1(_13434_),
    .A2(_13440_),
    .B1_N(_13438_),
    .Y(_13765_));
 sky130_fd_sc_hd__a31oi_4 _36333_ (.A1(_13759_),
    .A2(_13752_),
    .A3(_13757_),
    .B1(_13763_),
    .Y(_13766_));
 sky130_fd_sc_hd__a21o_1 _36334_ (.A1(_13752_),
    .A2(_13757_),
    .B1(_13759_),
    .X(_13767_));
 sky130_fd_sc_hd__nand2_1 _36335_ (.A(_13766_),
    .B(_13767_),
    .Y(_13768_));
 sky130_fd_sc_hd__nand3_4 _36336_ (.A(_13764_),
    .B(_13765_),
    .C(_13768_),
    .Y(_13769_));
 sky130_vsdinv _36337_ (.A(_13763_),
    .Y(_13770_));
 sky130_fd_sc_hd__o21ai_2 _36338_ (.A1(_13760_),
    .A2(_13762_),
    .B1(_13770_),
    .Y(_13771_));
 sky130_fd_sc_hd__nand2_1 _36339_ (.A(_13434_),
    .B(_13440_),
    .Y(_13772_));
 sky130_fd_sc_hd__nand2_1 _36340_ (.A(_13772_),
    .B(_13438_),
    .Y(_13773_));
 sky130_fd_sc_hd__nand3_1 _36341_ (.A(_13759_),
    .B(_13757_),
    .C(_13752_),
    .Y(_13774_));
 sky130_fd_sc_hd__nand3_2 _36342_ (.A(_13767_),
    .B(_13774_),
    .C(_13763_),
    .Y(_13775_));
 sky130_fd_sc_hd__nand3_4 _36343_ (.A(_13771_),
    .B(_13773_),
    .C(_13775_),
    .Y(_13776_));
 sky130_fd_sc_hd__nand2_4 _36344_ (.A(_19902_),
    .B(_11587_),
    .Y(_13777_));
 sky130_fd_sc_hd__nand2_4 _36345_ (.A(_19906_),
    .B(_20073_),
    .Y(_13778_));
 sky130_fd_sc_hd__nor2_8 _36346_ (.A(_13777_),
    .B(_13778_),
    .Y(_13779_));
 sky130_fd_sc_hd__nand2_2 _36347_ (.A(_19910_),
    .B(_11604_),
    .Y(_13780_));
 sky130_vsdinv _36348_ (.A(_13780_),
    .Y(_13781_));
 sky130_fd_sc_hd__nand2_1 _36349_ (.A(_13777_),
    .B(_13778_),
    .Y(_13782_));
 sky130_fd_sc_hd__nand3b_1 _36350_ (.A_N(_13779_),
    .B(_13781_),
    .C(_13782_),
    .Y(_13783_));
 sky130_fd_sc_hd__a22oi_1 _36351_ (.A1(_19903_),
    .A2(_20079_),
    .B1(_19907_),
    .B2(_11607_),
    .Y(_13784_));
 sky130_fd_sc_hd__o21ai_1 _36352_ (.A1(_13784_),
    .A2(_13779_),
    .B1(_13780_),
    .Y(_13785_));
 sky130_fd_sc_hd__nand2_2 _36353_ (.A(_13783_),
    .B(_13785_),
    .Y(_13786_));
 sky130_vsdinv _36354_ (.A(_13786_),
    .Y(_13787_));
 sky130_fd_sc_hd__nand2_2 _36355_ (.A(_10692_),
    .B(_09902_),
    .Y(_13788_));
 sky130_fd_sc_hd__a21o_1 _36356_ (.A1(_19897_),
    .A2(_20087_),
    .B1(_13788_),
    .X(_13789_));
 sky130_fd_sc_hd__nand2_2 _36357_ (.A(_10693_),
    .B(_20086_),
    .Y(_13790_));
 sky130_fd_sc_hd__a21o_1 _36358_ (.A1(_19894_),
    .A2(_11927_),
    .B1(_13790_),
    .X(_13791_));
 sky130_fd_sc_hd__nand2_2 _36359_ (.A(_19899_),
    .B(_11157_),
    .Y(_13792_));
 sky130_fd_sc_hd__nand3_4 _36360_ (.A(_13789_),
    .B(_13791_),
    .C(_13792_),
    .Y(_13793_));
 sky130_fd_sc_hd__nand3_2 _36361_ (.A(_19894_),
    .B(_19897_),
    .C(_13456_),
    .Y(_13794_));
 sky130_fd_sc_hd__nand2_4 _36362_ (.A(_13788_),
    .B(_13790_),
    .Y(_13795_));
 sky130_vsdinv _36363_ (.A(_13792_),
    .Y(_13796_));
 sky130_fd_sc_hd__o211ai_4 _36364_ (.A1(_12307_),
    .A2(_13794_),
    .B1(_13795_),
    .C1(_13796_),
    .Y(_13797_));
 sky130_fd_sc_hd__nand2_1 _36365_ (.A(_13793_),
    .B(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__a21oi_1 _36366_ (.A1(_13452_),
    .A2(_13450_),
    .B1(_13448_),
    .Y(_13799_));
 sky130_fd_sc_hd__nand2_2 _36367_ (.A(_13798_),
    .B(_13799_),
    .Y(_13800_));
 sky130_fd_sc_hd__o21bai_2 _36368_ (.A1(_13449_),
    .A2(_13454_),
    .B1_N(_13448_),
    .Y(_13801_));
 sky130_fd_sc_hd__nand3_4 _36369_ (.A(_13801_),
    .B(_13793_),
    .C(_13797_),
    .Y(_13802_));
 sky130_fd_sc_hd__and3_1 _36370_ (.A(_13787_),
    .B(_13800_),
    .C(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__a21oi_2 _36371_ (.A1(_13800_),
    .A2(_13802_),
    .B1(_13787_),
    .Y(_13804_));
 sky130_fd_sc_hd__o2bb2ai_4 _36372_ (.A1_N(_13769_),
    .A2_N(_13776_),
    .B1(_13803_),
    .B2(_13804_),
    .Y(_13805_));
 sky130_fd_sc_hd__a21o_1 _36373_ (.A1(_13800_),
    .A2(_13802_),
    .B1(_13786_),
    .X(_13806_));
 sky130_fd_sc_hd__nand3_1 _36374_ (.A(_13800_),
    .B(_13802_),
    .C(_13786_),
    .Y(_13807_));
 sky130_fd_sc_hd__nand2_2 _36375_ (.A(_13806_),
    .B(_13807_),
    .Y(_13808_));
 sky130_fd_sc_hd__nand3_4 _36376_ (.A(_13808_),
    .B(_13776_),
    .C(_13769_),
    .Y(_13809_));
 sky130_fd_sc_hd__nand2_1 _36377_ (.A(_13805_),
    .B(_13809_),
    .Y(_13810_));
 sky130_fd_sc_hd__nand2_1 _36378_ (.A(_13525_),
    .B(_13611_),
    .Y(_13811_));
 sky130_fd_sc_hd__nand2_1 _36379_ (.A(_13811_),
    .B(_13524_),
    .Y(_13812_));
 sky130_fd_sc_hd__nand2_4 _36380_ (.A(_13810_),
    .B(_13812_),
    .Y(_13813_));
 sky130_fd_sc_hd__a21oi_2 _36381_ (.A1(_13519_),
    .A2(_13521_),
    .B1(_13523_),
    .Y(_13814_));
 sky130_fd_sc_hd__o21ai_2 _36382_ (.A1(_13611_),
    .A2(_13814_),
    .B1(_13526_),
    .Y(_13815_));
 sky130_fd_sc_hd__nand3_4 _36383_ (.A(_13815_),
    .B(_13805_),
    .C(_13809_),
    .Y(_13816_));
 sky130_fd_sc_hd__a21boi_4 _36384_ (.A1(_13446_),
    .A2(_13483_),
    .B1_N(_13443_),
    .Y(_13817_));
 sky130_vsdinv _36385_ (.A(_13817_),
    .Y(_13818_));
 sky130_fd_sc_hd__a21oi_4 _36386_ (.A1(_13813_),
    .A2(_13816_),
    .B1(_13818_),
    .Y(_13819_));
 sky130_fd_sc_hd__nand3_2 _36387_ (.A(_13813_),
    .B(_13818_),
    .C(_13816_),
    .Y(_13820_));
 sky130_vsdinv _36388_ (.A(_13820_),
    .Y(_13821_));
 sky130_fd_sc_hd__a22oi_4 _36389_ (.A1(_09997_),
    .A2(_08008_),
    .B1(_09998_),
    .B2(net466),
    .Y(_13822_));
 sky130_fd_sc_hd__nor2_2 _36390_ (.A(_06155_),
    .B(net463),
    .Y(_13823_));
 sky130_fd_sc_hd__nand2_2 _36391_ (.A(_19844_),
    .B(_06312_),
    .Y(_13824_));
 sky130_vsdinv _36392_ (.A(_13824_),
    .Y(_13825_));
 sky130_fd_sc_hd__o21ai_1 _36393_ (.A1(_13822_),
    .A2(_13823_),
    .B1(_13825_),
    .Y(_13826_));
 sky130_vsdinv _36394_ (.A(_13826_),
    .Y(_13827_));
 sky130_fd_sc_hd__nor2_1 _36395_ (.A(_13822_),
    .B(_13823_),
    .Y(_13828_));
 sky130_fd_sc_hd__nand2_1 _36396_ (.A(_13828_),
    .B(_13824_),
    .Y(_13829_));
 sky130_vsdinv _36397_ (.A(_13829_),
    .Y(_13830_));
 sky130_fd_sc_hd__nand3_4 _36398_ (.A(_12487_),
    .B(_10972_),
    .C(_05820_),
    .Y(_13831_));
 sky130_fd_sc_hd__nor2_4 _36399_ (.A(_20153_),
    .B(_13831_),
    .Y(_13832_));
 sky130_fd_sc_hd__a22oi_4 _36400_ (.A1(_10972_),
    .A2(_10611_),
    .B1(_08242_),
    .B2(_10973_),
    .Y(_13833_));
 sky130_fd_sc_hd__nand2_4 _36401_ (.A(_19833_),
    .B(_05823_),
    .Y(_13834_));
 sky130_fd_sc_hd__o21ai_4 _36402_ (.A1(_13832_),
    .A2(_13833_),
    .B1(_13834_),
    .Y(_13835_));
 sky130_fd_sc_hd__nand2_2 _36403_ (.A(_12492_),
    .B(_05820_),
    .Y(_13836_));
 sky130_fd_sc_hd__buf_4 _36404_ (.A(_11778_),
    .X(_13837_));
 sky130_fd_sc_hd__nand3b_4 _36405_ (.A_N(_13836_),
    .B(_13837_),
    .C(_10446_),
    .Y(_13838_));
 sky130_fd_sc_hd__o21ai_4 _36406_ (.A1(_20153_),
    .A2(_11275_),
    .B1(_13836_),
    .Y(_13839_));
 sky130_vsdinv _36407_ (.A(_13834_),
    .Y(_13840_));
 sky130_fd_sc_hd__nand3_4 _36408_ (.A(_13838_),
    .B(_13839_),
    .C(_13840_),
    .Y(_13841_));
 sky130_fd_sc_hd__o21ai_4 _36409_ (.A1(_13571_),
    .A2(_13566_),
    .B1(_13569_),
    .Y(_13842_));
 sky130_fd_sc_hd__a21oi_4 _36410_ (.A1(_13835_),
    .A2(_13841_),
    .B1(_13842_),
    .Y(_13843_));
 sky130_fd_sc_hd__o21bai_2 _36411_ (.A1(_20153_),
    .A2(_13831_),
    .B1_N(_13834_),
    .Y(_13844_));
 sky130_fd_sc_hd__o211a_4 _36412_ (.A1(_13833_),
    .A2(_13844_),
    .B1(_13842_),
    .C1(_13835_),
    .X(_13845_));
 sky130_fd_sc_hd__o22ai_4 _36413_ (.A1(_13827_),
    .A2(_13830_),
    .B1(_13843_),
    .B2(_13845_),
    .Y(_13846_));
 sky130_fd_sc_hd__a21oi_2 _36414_ (.A1(_13582_),
    .A2(_13587_),
    .B1(_13576_),
    .Y(_13847_));
 sky130_fd_sc_hd__nor2_4 _36415_ (.A(_13833_),
    .B(_13844_),
    .Y(_13848_));
 sky130_fd_sc_hd__a21oi_2 _36416_ (.A1(_13838_),
    .A2(_13839_),
    .B1(_13840_),
    .Y(_13849_));
 sky130_fd_sc_hd__o21bai_4 _36417_ (.A1(_13848_),
    .A2(_13849_),
    .B1_N(_13842_),
    .Y(_13850_));
 sky130_fd_sc_hd__nand3_4 _36418_ (.A(_13835_),
    .B(_13842_),
    .C(_13841_),
    .Y(_13851_));
 sky130_fd_sc_hd__nand2_1 _36419_ (.A(_13828_),
    .B(_13825_),
    .Y(_13852_));
 sky130_fd_sc_hd__o21ai_1 _36420_ (.A1(_13822_),
    .A2(_13823_),
    .B1(_13824_),
    .Y(_13853_));
 sky130_fd_sc_hd__nand2_2 _36421_ (.A(_13852_),
    .B(_13853_),
    .Y(_13854_));
 sky130_fd_sc_hd__nand3_4 _36422_ (.A(_13850_),
    .B(_13851_),
    .C(_13854_),
    .Y(_13855_));
 sky130_fd_sc_hd__nand3_4 _36423_ (.A(_13846_),
    .B(_13847_),
    .C(_13855_),
    .Y(_13856_));
 sky130_fd_sc_hd__and2_1 _36424_ (.A(_13828_),
    .B(_13825_),
    .X(_13857_));
 sky130_vsdinv _36425_ (.A(_13853_),
    .Y(_13858_));
 sky130_fd_sc_hd__o22ai_4 _36426_ (.A1(_13857_),
    .A2(_13858_),
    .B1(_13843_),
    .B2(_13845_),
    .Y(_13859_));
 sky130_fd_sc_hd__o21ai_1 _36427_ (.A1(_13554_),
    .A2(_13558_),
    .B1(_13561_),
    .Y(_13860_));
 sky130_fd_sc_hd__o21ai_2 _36428_ (.A1(_13860_),
    .A2(_13574_),
    .B1(_13583_),
    .Y(_13861_));
 sky130_fd_sc_hd__nand2_2 _36429_ (.A(_13829_),
    .B(_13826_),
    .Y(_13862_));
 sky130_fd_sc_hd__nand3_2 _36430_ (.A(_13850_),
    .B(_13851_),
    .C(_13862_),
    .Y(_13863_));
 sky130_fd_sc_hd__nand3_4 _36431_ (.A(_13859_),
    .B(_13861_),
    .C(_13863_),
    .Y(_13864_));
 sky130_fd_sc_hd__nand2_1 _36432_ (.A(_13856_),
    .B(_13864_),
    .Y(_13865_));
 sky130_fd_sc_hd__nand2_2 _36433_ (.A(_19847_),
    .B(_06715_),
    .Y(_13866_));
 sky130_fd_sc_hd__a21o_1 _36434_ (.A1(_11363_),
    .A2(_12846_),
    .B1(_13866_),
    .X(_13867_));
 sky130_fd_sc_hd__nand2_1 _36435_ (.A(_10553_),
    .B(_20130_),
    .Y(_13868_));
 sky130_fd_sc_hd__a21o_1 _36436_ (.A1(_11366_),
    .A2(_20134_),
    .B1(_13868_),
    .X(_13869_));
 sky130_fd_sc_hd__nand2_2 _36437_ (.A(_19854_),
    .B(_07543_),
    .Y(_13870_));
 sky130_fd_sc_hd__nand3_4 _36438_ (.A(_13867_),
    .B(_13869_),
    .C(_13870_),
    .Y(_13871_));
 sky130_fd_sc_hd__nand3b_4 _36439_ (.A_N(_13866_),
    .B(_11010_),
    .C(_11093_),
    .Y(_13872_));
 sky130_vsdinv _36440_ (.A(_13870_),
    .Y(_13873_));
 sky130_fd_sc_hd__nand2_1 _36441_ (.A(_13866_),
    .B(_13868_),
    .Y(_13874_));
 sky130_fd_sc_hd__nand3_2 _36442_ (.A(_13872_),
    .B(_13873_),
    .C(_13874_),
    .Y(_13875_));
 sky130_fd_sc_hd__buf_4 _36443_ (.A(_13875_),
    .X(_13876_));
 sky130_fd_sc_hd__nor2_1 _36444_ (.A(_13556_),
    .B(_13554_),
    .Y(_13877_));
 sky130_fd_sc_hd__o2bb2ai_2 _36445_ (.A1_N(_13871_),
    .A2_N(_13876_),
    .B1(_13560_),
    .B2(_13877_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand2_4 _36446_ (.A(_13585_),
    .B(_13558_),
    .Y(_13879_));
 sky130_fd_sc_hd__nand3_4 _36447_ (.A(_13879_),
    .B(_13871_),
    .C(_13876_),
    .Y(_13880_));
 sky130_fd_sc_hd__a21oi_4 _36448_ (.A1(_13539_),
    .A2(_13538_),
    .B1(_13533_),
    .Y(_13881_));
 sky130_fd_sc_hd__a21oi_1 _36449_ (.A1(_13878_),
    .A2(_13880_),
    .B1(_13881_),
    .Y(_13882_));
 sky130_fd_sc_hd__a21oi_4 _36450_ (.A1(_13871_),
    .A2(_13876_),
    .B1(_13879_),
    .Y(_13883_));
 sky130_fd_sc_hd__nand2_2 _36451_ (.A(_13880_),
    .B(_13881_),
    .Y(_13884_));
 sky130_fd_sc_hd__nor2_1 _36452_ (.A(_13883_),
    .B(_13884_),
    .Y(_13885_));
 sky130_fd_sc_hd__nor2_1 _36453_ (.A(_13882_),
    .B(_13885_),
    .Y(_13886_));
 sky130_fd_sc_hd__nand2_2 _36454_ (.A(_13865_),
    .B(_13886_),
    .Y(_13887_));
 sky130_vsdinv _36455_ (.A(_13542_),
    .Y(_13888_));
 sky130_fd_sc_hd__nand2_4 _36456_ (.A(_13546_),
    .B(_13548_),
    .Y(_13889_));
 sky130_fd_sc_hd__nand2_1 _36457_ (.A(_13550_),
    .B(_13547_),
    .Y(_13890_));
 sky130_fd_sc_hd__o21ai_2 _36458_ (.A1(_13888_),
    .A2(_13889_),
    .B1(_13890_),
    .Y(_13891_));
 sky130_fd_sc_hd__o21ai_4 _36459_ (.A1(_13891_),
    .A2(_13591_),
    .B1(_13598_),
    .Y(_13892_));
 sky130_fd_sc_hd__nand2_1 _36460_ (.A(_13878_),
    .B(_13880_),
    .Y(_13893_));
 sky130_vsdinv _36461_ (.A(_13881_),
    .Y(_13894_));
 sky130_fd_sc_hd__o2bb2ai_4 _36462_ (.A1_N(_13893_),
    .A2_N(_13894_),
    .B1(_13883_),
    .B2(_13884_),
    .Y(_13895_));
 sky130_fd_sc_hd__nand3_4 _36463_ (.A(_13856_),
    .B(_13864_),
    .C(_13895_),
    .Y(_13896_));
 sky130_fd_sc_hd__nand3_4 _36464_ (.A(_13887_),
    .B(_13892_),
    .C(_13896_),
    .Y(_13897_));
 sky130_fd_sc_hd__a21oi_2 _36465_ (.A1(_13856_),
    .A2(_13864_),
    .B1(_13895_),
    .Y(_13898_));
 sky130_fd_sc_hd__o211a_1 _36466_ (.A1(_13882_),
    .A2(_13885_),
    .B1(_13864_),
    .C1(_13856_),
    .X(_13899_));
 sky130_fd_sc_hd__a21oi_2 _36467_ (.A1(_13596_),
    .A2(_13597_),
    .B1(_13594_),
    .Y(_13900_));
 sky130_fd_sc_hd__o21ai_4 _36468_ (.A1(_13898_),
    .A2(_13899_),
    .B1(_13900_),
    .Y(_13901_));
 sky130_fd_sc_hd__buf_4 _36469_ (.A(_08582_),
    .X(_13902_));
 sky130_fd_sc_hd__nand3_4 _36470_ (.A(_13902_),
    .B(_13497_),
    .C(_10694_),
    .Y(_13903_));
 sky130_fd_sc_hd__nor2_2 _36471_ (.A(_10691_),
    .B(_13903_),
    .Y(_13904_));
 sky130_fd_sc_hd__a22o_2 _36472_ (.A1(_11396_),
    .A2(_20124_),
    .B1(_12855_),
    .B2(_20119_),
    .X(_13905_));
 sky130_fd_sc_hd__nand2_4 _36473_ (.A(_19866_),
    .B(_08060_),
    .Y(_13906_));
 sky130_fd_sc_hd__nand3b_4 _36474_ (.A_N(_13904_),
    .B(_13905_),
    .C(_13906_),
    .Y(_13907_));
 sky130_fd_sc_hd__a21oi_2 _36475_ (.A1(_13498_),
    .A2(_13496_),
    .B1(_13494_),
    .Y(_13908_));
 sky130_fd_sc_hd__a22oi_4 _36476_ (.A1(_13902_),
    .A2(_09443_),
    .B1(_12447_),
    .B2(_07726_),
    .Y(_13909_));
 sky130_vsdinv _36477_ (.A(_13906_),
    .Y(_13910_));
 sky130_fd_sc_hd__o21ai_2 _36478_ (.A1(_13909_),
    .A2(_13904_),
    .B1(_13910_),
    .Y(_13911_));
 sky130_fd_sc_hd__nand3_4 _36479_ (.A(_13907_),
    .B(_13908_),
    .C(_13911_),
    .Y(_13912_));
 sky130_fd_sc_hd__nor2_2 _36480_ (.A(_13495_),
    .B(_13501_),
    .Y(_13913_));
 sky130_fd_sc_hd__o211ai_4 _36481_ (.A1(_10704_),
    .A2(_13903_),
    .B1(_13910_),
    .C1(_13905_),
    .Y(_13914_));
 sky130_fd_sc_hd__o21ai_2 _36482_ (.A1(_13909_),
    .A2(_13904_),
    .B1(_13906_),
    .Y(_13915_));
 sky130_fd_sc_hd__o211ai_4 _36483_ (.A1(_13494_),
    .A2(_13913_),
    .B1(_13914_),
    .C1(_13915_),
    .Y(_13916_));
 sky130_fd_sc_hd__nand2_2 _36484_ (.A(_12864_),
    .B(_11487_),
    .Y(_13917_));
 sky130_fd_sc_hd__nand3b_4 _36485_ (.A_N(_13917_),
    .B(_19875_),
    .C(_13758_),
    .Y(_13918_));
 sky130_fd_sc_hd__nand2_1 _36486_ (.A(_10936_),
    .B(_10343_),
    .Y(_13919_));
 sky130_fd_sc_hd__nand2_2 _36487_ (.A(_13917_),
    .B(_13919_),
    .Y(_13920_));
 sky130_fd_sc_hd__nand2_4 _36488_ (.A(_07479_),
    .B(_20105_),
    .Y(_13921_));
 sky130_fd_sc_hd__a21o_1 _36489_ (.A1(_13918_),
    .A2(_13920_),
    .B1(_13921_),
    .X(_13922_));
 sky130_fd_sc_hd__nand3_2 _36490_ (.A(_13918_),
    .B(_13921_),
    .C(_13920_),
    .Y(_13923_));
 sky130_fd_sc_hd__nand2_4 _36491_ (.A(_13922_),
    .B(_13923_),
    .Y(_13924_));
 sky130_fd_sc_hd__a21o_2 _36492_ (.A1(_13912_),
    .A2(_13916_),
    .B1(_13924_),
    .X(_13925_));
 sky130_fd_sc_hd__nand3_4 _36493_ (.A(_13924_),
    .B(_13916_),
    .C(_13912_),
    .Y(_13926_));
 sky130_fd_sc_hd__nand2_8 _36494_ (.A(_13889_),
    .B(_13542_),
    .Y(_13927_));
 sky130_fd_sc_hd__a21oi_4 _36495_ (.A1(_13925_),
    .A2(_13926_),
    .B1(_13927_),
    .Y(_13928_));
 sky130_vsdinv _36496_ (.A(_13916_),
    .Y(_13929_));
 sky130_fd_sc_hd__nand2_1 _36497_ (.A(_13924_),
    .B(_13912_),
    .Y(_13930_));
 sky130_fd_sc_hd__o211a_2 _36498_ (.A1(_13929_),
    .A2(_13930_),
    .B1(_13925_),
    .C1(_13927_),
    .X(_13931_));
 sky130_fd_sc_hd__nand2_1 _36499_ (.A(_13520_),
    .B(_13507_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand2_2 _36500_ (.A(_13932_),
    .B(_13503_),
    .Y(_13933_));
 sky130_vsdinv _36501_ (.A(_13933_),
    .Y(_13934_));
 sky130_fd_sc_hd__o21ai_2 _36502_ (.A1(_13928_),
    .A2(_13931_),
    .B1(_13934_),
    .Y(_13935_));
 sky130_vsdinv _36503_ (.A(_13935_),
    .Y(_13936_));
 sky130_fd_sc_hd__a21o_1 _36504_ (.A1(_13925_),
    .A2(_13926_),
    .B1(_13927_),
    .X(_13937_));
 sky130_fd_sc_hd__nand2_1 _36505_ (.A(_13937_),
    .B(_13933_),
    .Y(_13938_));
 sky130_fd_sc_hd__nor2_2 _36506_ (.A(_13931_),
    .B(_13938_),
    .Y(_13939_));
 sky130_fd_sc_hd__o2bb2ai_4 _36507_ (.A1_N(_13897_),
    .A2_N(_13901_),
    .B1(_13936_),
    .B2(_13939_),
    .Y(_13940_));
 sky130_fd_sc_hd__o21ai_1 _36508_ (.A1(_13928_),
    .A2(_13931_),
    .B1(_13933_),
    .Y(_13941_));
 sky130_fd_sc_hd__nand3_4 _36509_ (.A(_13927_),
    .B(_13925_),
    .C(_13926_),
    .Y(_13942_));
 sky130_fd_sc_hd__nand3_1 _36510_ (.A(_13937_),
    .B(_13942_),
    .C(_13934_),
    .Y(_13943_));
 sky130_fd_sc_hd__nand2_2 _36511_ (.A(_13941_),
    .B(_13943_),
    .Y(_13944_));
 sky130_fd_sc_hd__nand3_4 _36512_ (.A(_13901_),
    .B(_13897_),
    .C(_13944_),
    .Y(_13945_));
 sky130_fd_sc_hd__nor2_1 _36513_ (.A(_13611_),
    .B(_13814_),
    .Y(_13946_));
 sky130_fd_sc_hd__a21o_1 _36514_ (.A1(_13526_),
    .A2(_13946_),
    .B1(_13529_),
    .X(_13947_));
 sky130_fd_sc_hd__o21ai_4 _36515_ (.A1(_13602_),
    .A2(_13947_),
    .B1(_13610_),
    .Y(_13948_));
 sky130_fd_sc_hd__a21oi_4 _36516_ (.A1(_13940_),
    .A2(_13945_),
    .B1(_13948_),
    .Y(_13949_));
 sky130_fd_sc_hd__a22oi_1 _36517_ (.A1(_13612_),
    .A2(_13613_),
    .B1(_13607_),
    .B2(_13608_),
    .Y(_13950_));
 sky130_fd_sc_hd__o211a_1 _36518_ (.A1(_13605_),
    .A2(_13950_),
    .B1(_13945_),
    .C1(_13940_),
    .X(_13951_));
 sky130_fd_sc_hd__o22ai_4 _36519_ (.A1(_13819_),
    .A2(_13821_),
    .B1(_13949_),
    .B2(_13951_),
    .Y(_13952_));
 sky130_fd_sc_hd__a21o_2 _36520_ (.A1(_13940_),
    .A2(_13945_),
    .B1(_13948_),
    .X(_13953_));
 sky130_fd_sc_hd__nor2_2 _36521_ (.A(_13819_),
    .B(_13821_),
    .Y(_13954_));
 sky130_fd_sc_hd__nand3_4 _36522_ (.A(_13948_),
    .B(_13940_),
    .C(_13945_),
    .Y(_13955_));
 sky130_fd_sc_hd__nand3_2 _36523_ (.A(_13953_),
    .B(_13954_),
    .C(_13955_),
    .Y(_13956_));
 sky130_fd_sc_hd__nand3_4 _36524_ (.A(_13746_),
    .B(_13952_),
    .C(_13956_),
    .Y(_13957_));
 sky130_fd_sc_hd__a21oi_4 _36525_ (.A1(_13624_),
    .A2(_13627_),
    .B1(_13621_),
    .Y(_13958_));
 sky130_fd_sc_hd__o21ai_2 _36526_ (.A1(_13949_),
    .A2(_13951_),
    .B1(_13954_),
    .Y(_13959_));
 sky130_fd_sc_hd__a21o_1 _36527_ (.A1(_13813_),
    .A2(_13816_),
    .B1(_13818_),
    .X(_13960_));
 sky130_fd_sc_hd__nand2_2 _36528_ (.A(_13960_),
    .B(_13820_),
    .Y(_13961_));
 sky130_fd_sc_hd__nand3_2 _36529_ (.A(_13953_),
    .B(_13955_),
    .C(_13961_),
    .Y(_13962_));
 sky130_fd_sc_hd__nand3_4 _36530_ (.A(_13958_),
    .B(_13959_),
    .C(_13962_),
    .Y(_13963_));
 sky130_vsdinv _36531_ (.A(_13689_),
    .Y(_13964_));
 sky130_vsdinv _36532_ (.A(_13675_),
    .Y(_13965_));
 sky130_fd_sc_hd__nand2_2 _36533_ (.A(_13463_),
    .B(_13464_),
    .Y(_13966_));
 sky130_fd_sc_hd__a21o_1 _36534_ (.A1(_13468_),
    .A2(_13966_),
    .B1(_13465_),
    .X(_13967_));
 sky130_fd_sc_hd__o21ai_4 _36535_ (.A1(_07660_),
    .A2(_06840_),
    .B1(_18685_),
    .Y(_13968_));
 sky130_fd_sc_hd__and3_4 _36536_ (.A(_18685_),
    .B(_06659_),
    .C(_06110_),
    .X(_13969_));
 sky130_fd_sc_hd__o21ai_4 _36537_ (.A1(_13968_),
    .A2(_13969_),
    .B1(_13329_),
    .Y(_13970_));
 sky130_fd_sc_hd__o211a_4 _36538_ (.A1(_05722_),
    .A2(_05724_),
    .B1(_18685_),
    .C1(_19917_),
    .X(_13971_));
 sky130_fd_sc_hd__nand3_4 _36539_ (.A(net504),
    .B(_06095_),
    .C(_06657_),
    .Y(_13972_));
 sky130_fd_sc_hd__nand2_8 _36540_ (.A(_13971_),
    .B(_13972_),
    .Y(_13973_));
 sky130_fd_sc_hd__nand3_4 _36541_ (.A(_13967_),
    .B(_13970_),
    .C(_13973_),
    .Y(_13974_));
 sky130_fd_sc_hd__a21oi_4 _36542_ (.A1(_13468_),
    .A2(_13966_),
    .B1(_13465_),
    .Y(_13975_));
 sky130_fd_sc_hd__o21ai_4 _36543_ (.A1(_13968_),
    .A2(_13969_),
    .B1(_13324_),
    .Y(_13976_));
 sky130_fd_sc_hd__nand3b_4 _36544_ (.A_N(_13968_),
    .B(_13329_),
    .C(_13972_),
    .Y(_13977_));
 sky130_fd_sc_hd__nand3_4 _36545_ (.A(_13975_),
    .B(_13976_),
    .C(_13977_),
    .Y(_13978_));
 sky130_fd_sc_hd__a21o_2 _36546_ (.A1(_13325_),
    .A2(_13644_),
    .B1(_13640_),
    .X(_13979_));
 sky130_fd_sc_hd__a21oi_2 _36547_ (.A1(_13974_),
    .A2(_13978_),
    .B1(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__and3_1 _36548_ (.A(_13974_),
    .B(_13978_),
    .C(_13979_),
    .X(_13981_));
 sky130_fd_sc_hd__a21oi_4 _36549_ (.A1(_13475_),
    .A2(_13478_),
    .B1(_13461_),
    .Y(_13982_));
 sky130_fd_sc_hd__o21ai_4 _36550_ (.A1(_13980_),
    .A2(_13981_),
    .B1(_13982_),
    .Y(_13983_));
 sky130_fd_sc_hd__o2bb2ai_2 _36551_ (.A1_N(_13455_),
    .A2_N(_13473_),
    .B1(_13471_),
    .B2(_13458_),
    .Y(_13984_));
 sky130_fd_sc_hd__a21o_1 _36552_ (.A1(_13974_),
    .A2(_13978_),
    .B1(_13979_),
    .X(_13985_));
 sky130_fd_sc_hd__nand3_4 _36553_ (.A(_13974_),
    .B(_13978_),
    .C(_13979_),
    .Y(_13986_));
 sky130_fd_sc_hd__nand3_4 _36554_ (.A(_13984_),
    .B(_13985_),
    .C(_13986_),
    .Y(_13987_));
 sky130_fd_sc_hd__nand2_2 _36555_ (.A(_13653_),
    .B(_13656_),
    .Y(_13988_));
 sky130_fd_sc_hd__nand2_2 _36556_ (.A(_13988_),
    .B(_13649_),
    .Y(_13989_));
 sky130_fd_sc_hd__a21oi_4 _36557_ (.A1(_13983_),
    .A2(_13987_),
    .B1(_13989_),
    .Y(_13990_));
 sky130_vsdinv _36558_ (.A(_13649_),
    .Y(_13991_));
 sky130_fd_sc_hd__and2_1 _36559_ (.A(_13653_),
    .B(_13656_),
    .X(_13992_));
 sky130_fd_sc_hd__o211a_1 _36560_ (.A1(_13991_),
    .A2(_13992_),
    .B1(_13987_),
    .C1(_13983_),
    .X(_13993_));
 sky130_vsdinv _36561_ (.A(_13657_),
    .Y(_13994_));
 sky130_fd_sc_hd__nand2_1 _36562_ (.A(_13661_),
    .B(_13655_),
    .Y(_13995_));
 sky130_fd_sc_hd__a21oi_2 _36563_ (.A1(_13655_),
    .A2(_13657_),
    .B1(_13661_),
    .Y(_13996_));
 sky130_fd_sc_hd__o22ai_4 _36564_ (.A1(_13994_),
    .A2(_13995_),
    .B1(_13663_),
    .B2(_13996_),
    .Y(_13997_));
 sky130_fd_sc_hd__o21bai_4 _36565_ (.A1(_13990_),
    .A2(_13993_),
    .B1_N(_13997_),
    .Y(_13998_));
 sky130_fd_sc_hd__a21o_1 _36566_ (.A1(_13983_),
    .A2(_13987_),
    .B1(_13989_),
    .X(_13999_));
 sky130_fd_sc_hd__nand2_2 _36567_ (.A(_13985_),
    .B(_13986_),
    .Y(_14000_));
 sky130_fd_sc_hd__a22oi_4 _36568_ (.A1(_13649_),
    .A2(_13988_),
    .B1(_14000_),
    .B2(_13982_),
    .Y(_14001_));
 sky130_fd_sc_hd__nand2_2 _36569_ (.A(_14001_),
    .B(_13987_),
    .Y(_14002_));
 sky130_fd_sc_hd__nand3_4 _36570_ (.A(_13999_),
    .B(_14002_),
    .C(_13997_),
    .Y(_14003_));
 sky130_fd_sc_hd__a22oi_4 _36571_ (.A1(_13964_),
    .A2(_13965_),
    .B1(_13998_),
    .B2(_14003_),
    .Y(_14004_));
 sky130_fd_sc_hd__nand2_1 _36572_ (.A(_14002_),
    .B(_13997_),
    .Y(_14005_));
 sky130_fd_sc_hd__o211a_1 _36573_ (.A1(_13990_),
    .A2(_14005_),
    .B1(_13687_),
    .C1(_13998_),
    .X(_14006_));
 sky130_fd_sc_hd__o21a_2 _36574_ (.A1(_13489_),
    .A2(_13625_),
    .B1(_13488_),
    .X(_14007_));
 sky130_fd_sc_hd__o21ai_2 _36575_ (.A1(_14004_),
    .A2(_14006_),
    .B1(_14007_),
    .Y(_14008_));
 sky130_fd_sc_hd__buf_4 _36576_ (.A(_13677_),
    .X(_14009_));
 sky130_fd_sc_hd__a21o_1 _36577_ (.A1(_13998_),
    .A2(_14003_),
    .B1(_14009_),
    .X(_14010_));
 sky130_fd_sc_hd__nand3_4 _36578_ (.A(_13998_),
    .B(_13687_),
    .C(_14003_),
    .Y(_14011_));
 sky130_fd_sc_hd__o21ai_2 _36579_ (.A1(_13489_),
    .A2(_13625_),
    .B1(_13488_),
    .Y(_14012_));
 sky130_fd_sc_hd__nand3_4 _36580_ (.A(_14010_),
    .B(_14011_),
    .C(_14012_),
    .Y(_14013_));
 sky130_fd_sc_hd__buf_4 _36581_ (.A(_13686_),
    .X(_14014_));
 sky130_fd_sc_hd__a21bo_1 _36582_ (.A1(_14014_),
    .A2(_13668_),
    .B1_N(_13672_),
    .X(_14015_));
 sky130_fd_sc_hd__a21oi_4 _36583_ (.A1(_14008_),
    .A2(_14013_),
    .B1(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__clkbuf_4 _36584_ (.A(_14013_),
    .X(_14017_));
 sky130_fd_sc_hd__and3_2 _36585_ (.A(_14008_),
    .B(_14017_),
    .C(_14015_),
    .X(_14018_));
 sky130_fd_sc_hd__o2bb2ai_4 _36586_ (.A1_N(_13957_),
    .A2_N(_13963_),
    .B1(_14016_),
    .B2(_14018_),
    .Y(_14019_));
 sky130_fd_sc_hd__nand2_1 _36587_ (.A(_14010_),
    .B(_14011_),
    .Y(_14020_));
 sky130_fd_sc_hd__a21boi_4 _36588_ (.A1(_14020_),
    .A2(_14007_),
    .B1_N(_14015_),
    .Y(_14021_));
 sky130_fd_sc_hd__a21oi_4 _36589_ (.A1(_14017_),
    .A2(_14021_),
    .B1(_14016_),
    .Y(_14022_));
 sky130_fd_sc_hd__nand3_4 _36590_ (.A(_13963_),
    .B(_14022_),
    .C(_13957_),
    .Y(_14023_));
 sky130_fd_sc_hd__nand2_1 _36591_ (.A(_13637_),
    .B(_13701_),
    .Y(_14024_));
 sky130_fd_sc_hd__nand2_4 _36592_ (.A(_14024_),
    .B(_13630_),
    .Y(_14025_));
 sky130_fd_sc_hd__a21oi_4 _36593_ (.A1(_14019_),
    .A2(_14023_),
    .B1(_14025_),
    .Y(_14026_));
 sky130_vsdinv _36594_ (.A(_13957_),
    .Y(_14027_));
 sky130_fd_sc_hd__nand2_1 _36595_ (.A(_13963_),
    .B(_14022_),
    .Y(_14028_));
 sky130_fd_sc_hd__o211a_1 _36596_ (.A1(_14027_),
    .A2(_14028_),
    .B1(_14019_),
    .C1(_14025_),
    .X(_14029_));
 sky130_fd_sc_hd__o22ai_4 _36597_ (.A1(_13744_),
    .A2(_13745_),
    .B1(_14026_),
    .B2(_14029_),
    .Y(_14030_));
 sky130_fd_sc_hd__a21o_1 _36598_ (.A1(_14019_),
    .A2(_14023_),
    .B1(_14025_),
    .X(_14031_));
 sky130_fd_sc_hd__nand3_4 _36599_ (.A(_14025_),
    .B(_14019_),
    .C(_14023_),
    .Y(_14032_));
 sky130_fd_sc_hd__nor2_2 _36600_ (.A(_13744_),
    .B(_13745_),
    .Y(_14033_));
 sky130_fd_sc_hd__nand3_4 _36601_ (.A(_14031_),
    .B(_14032_),
    .C(_14033_),
    .Y(_14034_));
 sky130_fd_sc_hd__nand2_1 _36602_ (.A(_13708_),
    .B(_13718_),
    .Y(_14035_));
 sky130_fd_sc_hd__nand2_2 _36603_ (.A(_14035_),
    .B(_13703_),
    .Y(_14036_));
 sky130_fd_sc_hd__nand3_4 _36604_ (.A(_14030_),
    .B(_14034_),
    .C(_14036_),
    .Y(_14037_));
 sky130_fd_sc_hd__or2_2 _36605_ (.A(_13743_),
    .B(_13745_),
    .X(_14038_));
 sky130_fd_sc_hd__o21bai_2 _36606_ (.A1(_14026_),
    .A2(_14029_),
    .B1_N(_14038_),
    .Y(_14039_));
 sky130_fd_sc_hd__a21boi_4 _36607_ (.A1(_13708_),
    .A2(_13718_),
    .B1_N(_13703_),
    .Y(_14040_));
 sky130_fd_sc_hd__nand3_2 _36608_ (.A(_14031_),
    .B(_14032_),
    .C(_14038_),
    .Y(_14041_));
 sky130_fd_sc_hd__nand3_4 _36609_ (.A(_14039_),
    .B(_14040_),
    .C(_14041_),
    .Y(_14042_));
 sky130_fd_sc_hd__o2bb2ai_2 _36610_ (.A1_N(_14037_),
    .A2_N(_14042_),
    .B1(_13715_),
    .B2(_13710_),
    .Y(_14043_));
 sky130_fd_sc_hd__nand3_4 _36611_ (.A(_14042_),
    .B(_14037_),
    .C(_13717_),
    .Y(_14044_));
 sky130_fd_sc_hd__nand2_1 _36612_ (.A(_13720_),
    .B(_13405_),
    .Y(_14045_));
 sky130_fd_sc_hd__nand2_2 _36613_ (.A(_14045_),
    .B(_13724_),
    .Y(_14046_));
 sky130_fd_sc_hd__a21o_1 _36614_ (.A1(_14043_),
    .A2(_14044_),
    .B1(_14046_),
    .X(_14047_));
 sky130_fd_sc_hd__nand3_4 _36615_ (.A(_14043_),
    .B(_14046_),
    .C(_14044_),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_2 _36616_ (.A(_14047_),
    .B(_14048_),
    .Y(_14049_));
 sky130_fd_sc_hd__o2111ai_4 _36617_ (.A1(_13725_),
    .A2(_13729_),
    .B1(_13418_),
    .C1(_13734_),
    .D1(_13415_),
    .Y(_14050_));
 sky130_fd_sc_hd__nor2_4 _36618_ (.A(_14050_),
    .B(_13421_),
    .Y(_14051_));
 sky130_fd_sc_hd__and4_4 _36619_ (.A(_14051_),
    .B(_12052_),
    .C(_12053_),
    .D(_12422_),
    .X(_14052_));
 sky130_fd_sc_hd__a2bb2oi_2 _36620_ (.A1_N(_13725_),
    .A2_N(_13729_),
    .B1(_13734_),
    .B2(_13736_),
    .Y(_14053_));
 sky130_fd_sc_hd__o21ai_2 _36621_ (.A1(_14050_),
    .A2(_13423_),
    .B1(_14053_),
    .Y(_14054_));
 sky130_fd_sc_hd__a21oi_4 _36622_ (.A1(_12770_),
    .A2(_14051_),
    .B1(_14054_),
    .Y(_14055_));
 sky130_fd_sc_hd__a21boi_4 _36623_ (.A1(net409),
    .A2(_14052_),
    .B1_N(_14055_),
    .Y(_14056_));
 sky130_fd_sc_hd__or2_1 _36624_ (.A(_14049_),
    .B(_14056_),
    .X(_14057_));
 sky130_fd_sc_hd__nand2_1 _36625_ (.A(_14056_),
    .B(_14049_),
    .Y(_14058_));
 sky130_fd_sc_hd__and2_4 _36626_ (.A(_14057_),
    .B(_14058_),
    .X(_02659_));
 sky130_vsdinv _36627_ (.A(_14034_),
    .Y(_14059_));
 sky130_fd_sc_hd__nand2_1 _36628_ (.A(_14030_),
    .B(_14036_),
    .Y(_14060_));
 sky130_fd_sc_hd__o2bb2ai_1 _36629_ (.A1_N(_13717_),
    .A2_N(_14042_),
    .B1(_14059_),
    .B2(_14060_),
    .Y(_14061_));
 sky130_fd_sc_hd__a21boi_4 _36630_ (.A1(_13963_),
    .A2(_14022_),
    .B1_N(_13957_),
    .Y(_14062_));
 sky130_fd_sc_hd__nand2_2 _36631_ (.A(_13955_),
    .B(_13961_),
    .Y(_14063_));
 sky130_fd_sc_hd__o21ai_2 _36632_ (.A1(_13931_),
    .A2(_13938_),
    .B1(_13935_),
    .Y(_14064_));
 sky130_fd_sc_hd__a21oi_4 _36633_ (.A1(_13887_),
    .A2(_13896_),
    .B1(_13892_),
    .Y(_14065_));
 sky130_fd_sc_hd__o21ai_4 _36634_ (.A1(_14064_),
    .A2(_14065_),
    .B1(_13897_),
    .Y(_14066_));
 sky130_fd_sc_hd__a21oi_4 _36635_ (.A1(_13850_),
    .A2(_13862_),
    .B1(_13845_),
    .Y(_14067_));
 sky130_fd_sc_hd__nand2_2 _36636_ (.A(_09320_),
    .B(_07003_),
    .Y(_14068_));
 sky130_fd_sc_hd__a22oi_4 _36637_ (.A1(_10411_),
    .A2(_06151_),
    .B1(_19840_),
    .B2(_07004_),
    .Y(_14069_));
 sky130_fd_sc_hd__nand2_4 _36638_ (.A(_19835_),
    .B(_20138_),
    .Y(_14070_));
 sky130_fd_sc_hd__nand2_4 _36639_ (.A(_10989_),
    .B(_07503_),
    .Y(_14071_));
 sky130_fd_sc_hd__nor2_8 _36640_ (.A(_14070_),
    .B(_14071_),
    .Y(_14072_));
 sky130_fd_sc_hd__nor2_1 _36641_ (.A(_14069_),
    .B(_14072_),
    .Y(_14073_));
 sky130_fd_sc_hd__nor2_2 _36642_ (.A(_14068_),
    .B(_14073_),
    .Y(_14074_));
 sky130_fd_sc_hd__and2_1 _36643_ (.A(_14073_),
    .B(_14068_),
    .X(_14075_));
 sky130_fd_sc_hd__nand3_4 _36644_ (.A(_18693_),
    .B(_10575_),
    .C(_07033_),
    .Y(_14076_));
 sky130_fd_sc_hd__nor2_2 _36645_ (.A(_06148_),
    .B(_14076_),
    .Y(_14077_));
 sky130_fd_sc_hd__a22oi_4 _36646_ (.A1(_11783_),
    .A2(_05835_),
    .B1(_06672_),
    .B2(_11778_),
    .Y(_14078_));
 sky130_fd_sc_hd__o22ai_4 _36647_ (.A1(_10403_),
    .A2(_05813_),
    .B1(_14077_),
    .B2(_14078_),
    .Y(_14079_));
 sky130_fd_sc_hd__nand2_1 _36648_ (.A(_19828_),
    .B(_05822_),
    .Y(_14080_));
 sky130_fd_sc_hd__nand3b_4 _36649_ (.A_N(_14080_),
    .B(_12487_),
    .C(_06672_),
    .Y(_14081_));
 sky130_fd_sc_hd__o21ai_2 _36650_ (.A1(_10611_),
    .A2(_10968_),
    .B1(_14080_),
    .Y(_14082_));
 sky130_fd_sc_hd__nand2_4 _36651_ (.A(_10577_),
    .B(_20142_),
    .Y(_14083_));
 sky130_vsdinv _36652_ (.A(_14083_),
    .Y(_14084_));
 sky130_fd_sc_hd__nand3_4 _36653_ (.A(_14081_),
    .B(_14082_),
    .C(_14084_),
    .Y(_14085_));
 sky130_fd_sc_hd__o22ai_4 _36654_ (.A1(_20153_),
    .A2(_13831_),
    .B1(_13834_),
    .B2(_13833_),
    .Y(_14086_));
 sky130_fd_sc_hd__a21oi_4 _36655_ (.A1(_14079_),
    .A2(_14085_),
    .B1(_14086_),
    .Y(_14087_));
 sky130_fd_sc_hd__o21ai_1 _36656_ (.A1(net454),
    .A2(_14076_),
    .B1(_14084_),
    .Y(_14088_));
 sky130_fd_sc_hd__o211a_2 _36657_ (.A1(_14078_),
    .A2(_14088_),
    .B1(_14086_),
    .C1(_14079_),
    .X(_14089_));
 sky130_fd_sc_hd__o22ai_4 _36658_ (.A1(_14074_),
    .A2(_14075_),
    .B1(_14087_),
    .B2(_14089_),
    .Y(_14090_));
 sky130_fd_sc_hd__nand2_1 _36659_ (.A(_14079_),
    .B(_14085_),
    .Y(_14091_));
 sky130_fd_sc_hd__a21oi_4 _36660_ (.A1(_13839_),
    .A2(_13840_),
    .B1(_13832_),
    .Y(_14092_));
 sky130_fd_sc_hd__nand2_4 _36661_ (.A(_14091_),
    .B(_14092_),
    .Y(_14093_));
 sky130_fd_sc_hd__nand3_4 _36662_ (.A(_14079_),
    .B(_14086_),
    .C(_14085_),
    .Y(_14094_));
 sky130_fd_sc_hd__a21o_1 _36663_ (.A1(_14070_),
    .A2(_14071_),
    .B1(_14068_),
    .X(_14095_));
 sky130_fd_sc_hd__o21ai_2 _36664_ (.A1(_14069_),
    .A2(_14072_),
    .B1(_14068_),
    .Y(_14096_));
 sky130_fd_sc_hd__o21ai_4 _36665_ (.A1(_14072_),
    .A2(_14095_),
    .B1(_14096_),
    .Y(_14097_));
 sky130_fd_sc_hd__nand3_4 _36666_ (.A(_14093_),
    .B(_14094_),
    .C(_14097_),
    .Y(_14098_));
 sky130_fd_sc_hd__nand3_4 _36667_ (.A(_14067_),
    .B(_14090_),
    .C(_14098_),
    .Y(_14099_));
 sky130_fd_sc_hd__o21ai_2 _36668_ (.A1(_14087_),
    .A2(_14089_),
    .B1(_14097_),
    .Y(_14100_));
 sky130_fd_sc_hd__nand2_1 _36669_ (.A(_13835_),
    .B(_13842_),
    .Y(_14101_));
 sky130_fd_sc_hd__o22ai_4 _36670_ (.A1(_13848_),
    .A2(_14101_),
    .B1(_13854_),
    .B2(_13843_),
    .Y(_14102_));
 sky130_fd_sc_hd__o21a_1 _36671_ (.A1(_14072_),
    .A2(_14095_),
    .B1(_14096_),
    .X(_14103_));
 sky130_fd_sc_hd__nand3_2 _36672_ (.A(_14093_),
    .B(_14094_),
    .C(_14103_),
    .Y(_14104_));
 sky130_fd_sc_hd__nand3_4 _36673_ (.A(_14100_),
    .B(_14102_),
    .C(_14104_),
    .Y(_14105_));
 sky130_fd_sc_hd__nand2_1 _36674_ (.A(_14099_),
    .B(_14105_),
    .Y(_14106_));
 sky130_fd_sc_hd__nand2_2 _36675_ (.A(_10383_),
    .B(_06714_),
    .Y(_14107_));
 sky130_fd_sc_hd__nand3b_4 _36676_ (.A_N(_14107_),
    .B(_11363_),
    .C(_10350_),
    .Y(_14108_));
 sky130_fd_sc_hd__nand2_2 _36677_ (.A(_19854_),
    .B(_10694_),
    .Y(_14109_));
 sky130_vsdinv _36678_ (.A(_14109_),
    .Y(_14110_));
 sky130_fd_sc_hd__a22o_1 _36679_ (.A1(_11366_),
    .A2(_12846_),
    .B1(_12818_),
    .B2(_10350_),
    .X(_14111_));
 sky130_fd_sc_hd__nand3_4 _36680_ (.A(_14108_),
    .B(_14110_),
    .C(_14111_),
    .Y(_14112_));
 sky130_fd_sc_hd__a21o_1 _36681_ (.A1(_11363_),
    .A2(_10350_),
    .B1(_14107_),
    .X(_14113_));
 sky130_fd_sc_hd__nand3_4 _36682_ (.A(_14107_),
    .B(_19852_),
    .C(_20127_),
    .Y(_14114_));
 sky130_fd_sc_hd__nand3_4 _36683_ (.A(_14113_),
    .B(_14109_),
    .C(_14114_),
    .Y(_14115_));
 sky130_fd_sc_hd__o22ai_4 _36684_ (.A1(_06155_),
    .A2(_10988_),
    .B1(_13824_),
    .B2(_13822_),
    .Y(_14116_));
 sky130_fd_sc_hd__a21oi_4 _36685_ (.A1(_14112_),
    .A2(_14115_),
    .B1(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__a21oi_4 _36686_ (.A1(_13872_),
    .A2(_13876_),
    .B1(_14117_),
    .Y(_14118_));
 sky130_fd_sc_hd__nand3_4 _36687_ (.A(_14112_),
    .B(_14115_),
    .C(_14116_),
    .Y(_14119_));
 sky130_fd_sc_hd__nor2_1 _36688_ (.A(_13825_),
    .B(_13823_),
    .Y(_14120_));
 sky130_fd_sc_hd__o2bb2ai_2 _36689_ (.A1_N(_14115_),
    .A2_N(_14112_),
    .B1(_13822_),
    .B2(_14120_),
    .Y(_14121_));
 sky130_fd_sc_hd__nand2_1 _36690_ (.A(_13876_),
    .B(_13872_),
    .Y(_14122_));
 sky130_fd_sc_hd__a21oi_4 _36691_ (.A1(_14121_),
    .A2(_14119_),
    .B1(_14122_),
    .Y(_14123_));
 sky130_fd_sc_hd__a21oi_4 _36692_ (.A1(_14118_),
    .A2(_14119_),
    .B1(_14123_),
    .Y(_14124_));
 sky130_fd_sc_hd__nand2_1 _36693_ (.A(_14106_),
    .B(_14124_),
    .Y(_14125_));
 sky130_fd_sc_hd__a22oi_4 _36694_ (.A1(_13583_),
    .A2(_13588_),
    .B1(_13846_),
    .B2(_13855_),
    .Y(_14126_));
 sky130_fd_sc_hd__a21oi_4 _36695_ (.A1(_13856_),
    .A2(_13895_),
    .B1(_14126_),
    .Y(_14127_));
 sky130_fd_sc_hd__a21o_1 _36696_ (.A1(_14118_),
    .A2(_14119_),
    .B1(_14123_),
    .X(_14128_));
 sky130_fd_sc_hd__nand3_2 _36697_ (.A(_14128_),
    .B(_14099_),
    .C(_14105_),
    .Y(_14129_));
 sky130_fd_sc_hd__nand3_4 _36698_ (.A(_14125_),
    .B(_14127_),
    .C(_14129_),
    .Y(_14130_));
 sky130_fd_sc_hd__nand2_2 _36699_ (.A(_14106_),
    .B(_14128_),
    .Y(_14131_));
 sky130_fd_sc_hd__nand2_1 _36700_ (.A(_13856_),
    .B(_13895_),
    .Y(_14132_));
 sky130_fd_sc_hd__nand2_2 _36701_ (.A(_14132_),
    .B(_13864_),
    .Y(_14133_));
 sky130_fd_sc_hd__nand3_4 _36702_ (.A(_14099_),
    .B(_14105_),
    .C(_14124_),
    .Y(_14134_));
 sky130_fd_sc_hd__nand3_4 _36703_ (.A(_14131_),
    .B(_14133_),
    .C(_14134_),
    .Y(_14135_));
 sky130_fd_sc_hd__a31oi_4 _36704_ (.A1(_13879_),
    .A2(_13871_),
    .A3(_13876_),
    .B1(_13894_),
    .Y(_14136_));
 sky130_fd_sc_hd__o22ai_4 _36705_ (.A1(_10691_),
    .A2(_13903_),
    .B1(_13906_),
    .B2(_13909_),
    .Y(_14137_));
 sky130_fd_sc_hd__a22oi_4 _36706_ (.A1(_10440_),
    .A2(_12059_),
    .B1(_13497_),
    .B2(_10113_),
    .Y(_14138_));
 sky130_fd_sc_hd__nand3_4 _36707_ (.A(_10440_),
    .B(_10620_),
    .C(_12059_),
    .Y(_14139_));
 sky130_fd_sc_hd__nor2_2 _36708_ (.A(_12073_),
    .B(_14139_),
    .Y(_14140_));
 sky130_fd_sc_hd__nand2_4 _36709_ (.A(_19866_),
    .B(_07723_),
    .Y(_14141_));
 sky130_vsdinv _36710_ (.A(_14141_),
    .Y(_14142_));
 sky130_fd_sc_hd__o21ai_2 _36711_ (.A1(_14138_),
    .A2(_14140_),
    .B1(_14142_),
    .Y(_14143_));
 sky130_fd_sc_hd__a22o_2 _36712_ (.A1(_19859_),
    .A2(_11061_),
    .B1(_10926_),
    .B2(_11062_),
    .X(_14144_));
 sky130_fd_sc_hd__o211ai_4 _36713_ (.A1(_11074_),
    .A2(_14139_),
    .B1(_14141_),
    .C1(_14144_),
    .Y(_14145_));
 sky130_fd_sc_hd__nand3b_4 _36714_ (.A_N(_14137_),
    .B(_14143_),
    .C(_14145_),
    .Y(_14146_));
 sky130_fd_sc_hd__o21ai_2 _36715_ (.A1(_14138_),
    .A2(_14140_),
    .B1(_14141_),
    .Y(_14147_));
 sky130_fd_sc_hd__o211ai_4 _36716_ (.A1(_12073_),
    .A2(_14139_),
    .B1(_14142_),
    .C1(_14144_),
    .Y(_14148_));
 sky130_fd_sc_hd__nand3_4 _36717_ (.A(_14147_),
    .B(_14137_),
    .C(_14148_),
    .Y(_14149_));
 sky130_fd_sc_hd__a22oi_4 _36718_ (.A1(_12864_),
    .A2(_11723_),
    .B1(_11871_),
    .B2(_10716_),
    .Y(_14150_));
 sky130_fd_sc_hd__nand2_1 _36719_ (.A(_10628_),
    .B(_20107_),
    .Y(_14151_));
 sky130_fd_sc_hd__nand2_1 _36720_ (.A(_10944_),
    .B(_08450_),
    .Y(_14152_));
 sky130_fd_sc_hd__nor2_2 _36721_ (.A(_14151_),
    .B(_14152_),
    .Y(_14153_));
 sky130_fd_sc_hd__a211o_1 _36722_ (.A1(net457),
    .A2(_20103_),
    .B1(_14150_),
    .C1(_14153_),
    .X(_14154_));
 sky130_fd_sc_hd__clkbuf_4 _36723_ (.A(_14150_),
    .X(_14155_));
 sky130_fd_sc_hd__buf_2 _36724_ (.A(_14153_),
    .X(_14156_));
 sky130_fd_sc_hd__nand2_2 _36725_ (.A(_07479_),
    .B(_10811_),
    .Y(_14157_));
 sky130_vsdinv _36726_ (.A(_14157_),
    .Y(_14158_));
 sky130_fd_sc_hd__o21ai_1 _36727_ (.A1(_14155_),
    .A2(_14156_),
    .B1(_14158_),
    .Y(_14159_));
 sky130_fd_sc_hd__nand2_2 _36728_ (.A(_14154_),
    .B(_14159_),
    .Y(_14160_));
 sky130_fd_sc_hd__a21oi_4 _36729_ (.A1(_14146_),
    .A2(_14149_),
    .B1(_14160_),
    .Y(_14161_));
 sky130_fd_sc_hd__o21a_1 _36730_ (.A1(_14155_),
    .A2(_14156_),
    .B1(_14158_),
    .X(_14162_));
 sky130_fd_sc_hd__nor3_4 _36731_ (.A(_14158_),
    .B(_14155_),
    .C(_14156_),
    .Y(_14163_));
 sky130_fd_sc_hd__o211a_2 _36732_ (.A1(_14162_),
    .A2(_14163_),
    .B1(_14149_),
    .C1(_14146_),
    .X(_14164_));
 sky130_fd_sc_hd__o22ai_4 _36733_ (.A1(_13883_),
    .A2(_14136_),
    .B1(_14161_),
    .B2(_14164_),
    .Y(_14165_));
 sky130_fd_sc_hd__nand2_1 _36734_ (.A(_14146_),
    .B(_14149_),
    .Y(_14166_));
 sky130_fd_sc_hd__nor2_1 _36735_ (.A(_14163_),
    .B(_14162_),
    .Y(_14167_));
 sky130_fd_sc_hd__nand2_2 _36736_ (.A(_14166_),
    .B(_14167_),
    .Y(_14168_));
 sky130_fd_sc_hd__o21ai_4 _36737_ (.A1(_13881_),
    .A2(_13883_),
    .B1(_13880_),
    .Y(_14169_));
 sky130_fd_sc_hd__nand3_4 _36738_ (.A(_14160_),
    .B(_14146_),
    .C(_14149_),
    .Y(_14170_));
 sky130_fd_sc_hd__nand3_4 _36739_ (.A(_14168_),
    .B(_14169_),
    .C(_14170_),
    .Y(_14171_));
 sky130_fd_sc_hd__nand2_2 _36740_ (.A(_13930_),
    .B(_13916_),
    .Y(_14172_));
 sky130_fd_sc_hd__a21oi_4 _36741_ (.A1(_14165_),
    .A2(_14171_),
    .B1(_14172_),
    .Y(_14173_));
 sky130_vsdinv _36742_ (.A(_14171_),
    .Y(_14174_));
 sky130_fd_sc_hd__nand2_2 _36743_ (.A(_14165_),
    .B(_14172_),
    .Y(_14175_));
 sky130_fd_sc_hd__nor2_2 _36744_ (.A(_14174_),
    .B(_14175_),
    .Y(_14176_));
 sky130_fd_sc_hd__o2bb2ai_4 _36745_ (.A1_N(_14130_),
    .A2_N(_14135_),
    .B1(_14173_),
    .B2(_14176_),
    .Y(_14177_));
 sky130_fd_sc_hd__nand2_1 _36746_ (.A(_14168_),
    .B(_14170_),
    .Y(_14178_));
 sky130_fd_sc_hd__nand2_2 _36747_ (.A(_13884_),
    .B(_13878_),
    .Y(_14179_));
 sky130_fd_sc_hd__a21boi_4 _36748_ (.A1(_14178_),
    .A2(_14179_),
    .B1_N(_14172_),
    .Y(_14180_));
 sky130_fd_sc_hd__a21oi_4 _36749_ (.A1(_14171_),
    .A2(_14180_),
    .B1(_14173_),
    .Y(_14181_));
 sky130_fd_sc_hd__nand3_4 _36750_ (.A(_14135_),
    .B(_14130_),
    .C(_14181_),
    .Y(_14182_));
 sky130_fd_sc_hd__nand3_4 _36751_ (.A(_14066_),
    .B(_14177_),
    .C(_14182_),
    .Y(_14183_));
 sky130_fd_sc_hd__a21boi_4 _36752_ (.A1(_13901_),
    .A2(_13944_),
    .B1_N(_13897_),
    .Y(_14184_));
 sky130_fd_sc_hd__nand2_1 _36753_ (.A(_14135_),
    .B(_14130_),
    .Y(_14185_));
 sky130_fd_sc_hd__nand2_1 _36754_ (.A(_14185_),
    .B(_14181_),
    .Y(_14186_));
 sky130_fd_sc_hd__nand3b_2 _36755_ (.A_N(_14181_),
    .B(_14130_),
    .C(_14135_),
    .Y(_14187_));
 sky130_fd_sc_hd__nand3_4 _36756_ (.A(_14184_),
    .B(_14186_),
    .C(_14187_),
    .Y(_14188_));
 sky130_fd_sc_hd__a31oi_4 _36757_ (.A1(_13927_),
    .A2(_13925_),
    .A3(_13926_),
    .B1(_13933_),
    .Y(_14189_));
 sky130_fd_sc_hd__a22oi_4 _36758_ (.A1(_11463_),
    .A2(_09493_),
    .B1(_11455_),
    .B2(_12109_),
    .Y(_14190_));
 sky130_fd_sc_hd__nand3_4 _36759_ (.A(_11092_),
    .B(_12576_),
    .C(_12103_),
    .Y(_14191_));
 sky130_fd_sc_hd__nor2_8 _36760_ (.A(_11549_),
    .B(_14191_),
    .Y(_14192_));
 sky130_fd_sc_hd__nand2_4 _36761_ (.A(_19890_),
    .B(_11210_),
    .Y(_14193_));
 sky130_fd_sc_hd__o21ai_2 _36762_ (.A1(_14190_),
    .A2(_14192_),
    .B1(_14193_),
    .Y(_14194_));
 sky130_vsdinv _36763_ (.A(_14193_),
    .Y(_14195_));
 sky130_fd_sc_hd__a22o_2 _36764_ (.A1(_11463_),
    .A2(_11205_),
    .B1(_11455_),
    .B2(_12109_),
    .X(_14196_));
 sky130_fd_sc_hd__o211ai_4 _36765_ (.A1(_11563_),
    .A2(_14191_),
    .B1(_14195_),
    .C1(_14196_),
    .Y(_14197_));
 sky130_fd_sc_hd__a22oi_4 _36766_ (.A1(_19871_),
    .A2(_11492_),
    .B1(_19875_),
    .B2(_13758_),
    .Y(_14198_));
 sky130_fd_sc_hd__o21ai_4 _36767_ (.A1(_13921_),
    .A2(_14198_),
    .B1(_13918_),
    .Y(_14199_));
 sky130_fd_sc_hd__nand3_4 _36768_ (.A(_14194_),
    .B(_14197_),
    .C(_14199_),
    .Y(_14200_));
 sky130_fd_sc_hd__o21ai_4 _36769_ (.A1(_14190_),
    .A2(_14192_),
    .B1(_14195_),
    .Y(_14201_));
 sky130_fd_sc_hd__o21ai_2 _36770_ (.A1(_13917_),
    .A2(_13919_),
    .B1(_13921_),
    .Y(_14202_));
 sky130_fd_sc_hd__nand2_4 _36771_ (.A(_14202_),
    .B(_13920_),
    .Y(_14203_));
 sky130_fd_sc_hd__o211ai_4 _36772_ (.A1(_11557_),
    .A2(_14191_),
    .B1(_14193_),
    .C1(_14196_),
    .Y(_14204_));
 sky130_fd_sc_hd__nand3_4 _36773_ (.A(_14201_),
    .B(_14203_),
    .C(_14204_),
    .Y(_14205_));
 sky130_fd_sc_hd__nand2_2 _36774_ (.A(_13756_),
    .B(_13753_),
    .Y(_14206_));
 sky130_fd_sc_hd__a21oi_2 _36775_ (.A1(_14200_),
    .A2(_14205_),
    .B1(_14206_),
    .Y(_14207_));
 sky130_fd_sc_hd__and3_1 _36776_ (.A(_14200_),
    .B(_14205_),
    .C(_14206_),
    .X(_14208_));
 sky130_fd_sc_hd__o22ai_4 _36777_ (.A1(_13760_),
    .A2(_13766_),
    .B1(_14207_),
    .B2(_14208_),
    .Y(_14209_));
 sky130_fd_sc_hd__nor2_4 _36778_ (.A(_13760_),
    .B(_13766_),
    .Y(_14210_));
 sky130_fd_sc_hd__a21o_1 _36779_ (.A1(_14200_),
    .A2(_14205_),
    .B1(_14206_),
    .X(_14211_));
 sky130_fd_sc_hd__a32oi_4 _36780_ (.A1(_14201_),
    .A2(_14203_),
    .A3(_14204_),
    .B1(_13753_),
    .B2(_13757_),
    .Y(_14212_));
 sky130_fd_sc_hd__nand2_2 _36781_ (.A(_14212_),
    .B(_14200_),
    .Y(_14213_));
 sky130_fd_sc_hd__nand3_4 _36782_ (.A(_14210_),
    .B(_14211_),
    .C(_14213_),
    .Y(_14214_));
 sky130_fd_sc_hd__a22oi_4 _36783_ (.A1(_19894_),
    .A2(_10262_),
    .B1(_19897_),
    .B2(_12298_),
    .Y(_14215_));
 sky130_fd_sc_hd__nand3_4 _36784_ (.A(_11486_),
    .B(_07115_),
    .C(_09899_),
    .Y(_14216_));
 sky130_fd_sc_hd__nor2_4 _36785_ (.A(_09775_),
    .B(_14216_),
    .Y(_14217_));
 sky130_fd_sc_hd__nand2_2 _36786_ (.A(_19899_),
    .B(_10256_),
    .Y(_14218_));
 sky130_fd_sc_hd__o21ai_4 _36787_ (.A1(_14215_),
    .A2(_14217_),
    .B1(_14218_),
    .Y(_14219_));
 sky130_vsdinv _36788_ (.A(_14218_),
    .Y(_14220_));
 sky130_fd_sc_hd__a22o_2 _36789_ (.A1(_10692_),
    .A2(_20086_),
    .B1(_10693_),
    .B2(_20082_),
    .X(_14221_));
 sky130_fd_sc_hd__o211ai_4 _36790_ (.A1(_10763_),
    .A2(_14216_),
    .B1(_14220_),
    .C1(_14221_),
    .Y(_14222_));
 sky130_fd_sc_hd__nor2_2 _36791_ (.A(_13788_),
    .B(_13790_),
    .Y(_14223_));
 sky130_fd_sc_hd__a21o_2 _36792_ (.A1(_13796_),
    .A2(_13795_),
    .B1(_14223_),
    .X(_14224_));
 sky130_fd_sc_hd__a21oi_4 _36793_ (.A1(_14219_),
    .A2(_14222_),
    .B1(_14224_),
    .Y(_14225_));
 sky130_fd_sc_hd__a21oi_4 _36794_ (.A1(_13796_),
    .A2(_13795_),
    .B1(_14223_),
    .Y(_14226_));
 sky130_fd_sc_hd__nand2_1 _36795_ (.A(_14219_),
    .B(_14222_),
    .Y(_14227_));
 sky130_fd_sc_hd__nor2_2 _36796_ (.A(_14226_),
    .B(_14227_),
    .Y(_14228_));
 sky130_fd_sc_hd__a22oi_4 _36797_ (.A1(_10337_),
    .A2(_11174_),
    .B1(_10338_),
    .B2(_10778_),
    .Y(_14229_));
 sky130_fd_sc_hd__nand2_4 _36798_ (.A(_19902_),
    .B(_11173_),
    .Y(_14230_));
 sky130_fd_sc_hd__nand2_4 _36799_ (.A(_06107_),
    .B(_10777_),
    .Y(_14231_));
 sky130_fd_sc_hd__nor2_8 _36800_ (.A(_14230_),
    .B(_14231_),
    .Y(_14232_));
 sky130_fd_sc_hd__a211o_1 _36801_ (.A1(_18687_),
    .A2(_19910_),
    .B1(_14229_),
    .C1(_14232_),
    .X(_14233_));
 sky130_fd_sc_hd__nand2_8 _36802_ (.A(net504),
    .B(_05952_),
    .Y(_14234_));
 sky130_vsdinv _36803_ (.A(_14234_),
    .Y(_14235_));
 sky130_fd_sc_hd__o21ai_1 _36804_ (.A1(_14229_),
    .A2(_14232_),
    .B1(_14235_),
    .Y(_14236_));
 sky130_fd_sc_hd__nand2_1 _36805_ (.A(_14233_),
    .B(_14236_),
    .Y(_14237_));
 sky130_fd_sc_hd__o21ai_2 _36806_ (.A1(_14225_),
    .A2(_14228_),
    .B1(_14237_),
    .Y(_14238_));
 sky130_fd_sc_hd__nand2_2 _36807_ (.A(_14227_),
    .B(_14226_),
    .Y(_14239_));
 sky130_fd_sc_hd__nand3_4 _36808_ (.A(_14224_),
    .B(_14219_),
    .C(_14222_),
    .Y(_14240_));
 sky130_fd_sc_hd__nor3_4 _36809_ (.A(_14235_),
    .B(_14229_),
    .C(_14232_),
    .Y(_14241_));
 sky130_fd_sc_hd__o21a_2 _36810_ (.A1(_14229_),
    .A2(_14232_),
    .B1(_14235_),
    .X(_14242_));
 sky130_fd_sc_hd__nor2_8 _36811_ (.A(_14241_),
    .B(_14242_),
    .Y(_14243_));
 sky130_fd_sc_hd__nand3_4 _36812_ (.A(_14239_),
    .B(_14240_),
    .C(_14243_),
    .Y(_14244_));
 sky130_fd_sc_hd__nand2_4 _36813_ (.A(_14238_),
    .B(_14244_),
    .Y(_14245_));
 sky130_fd_sc_hd__a21oi_4 _36814_ (.A1(_14209_),
    .A2(_14214_),
    .B1(_14245_),
    .Y(_14246_));
 sky130_fd_sc_hd__a21oi_2 _36815_ (.A1(_14239_),
    .A2(_14240_),
    .B1(_14243_),
    .Y(_14247_));
 sky130_vsdinv _36816_ (.A(_14244_),
    .Y(_14248_));
 sky130_fd_sc_hd__o211a_1 _36817_ (.A1(_14247_),
    .A2(_14248_),
    .B1(_14214_),
    .C1(_14209_),
    .X(_14249_));
 sky130_fd_sc_hd__o22ai_4 _36818_ (.A1(_13928_),
    .A2(_14189_),
    .B1(_14246_),
    .B2(_14249_),
    .Y(_14250_));
 sky130_fd_sc_hd__o21ai_4 _36819_ (.A1(_13934_),
    .A2(_13928_),
    .B1(_13942_),
    .Y(_14251_));
 sky130_fd_sc_hd__a21o_1 _36820_ (.A1(_14209_),
    .A2(_14214_),
    .B1(_14245_),
    .X(_14252_));
 sky130_fd_sc_hd__nand3_4 _36821_ (.A(_14245_),
    .B(_14209_),
    .C(_14214_),
    .Y(_14253_));
 sky130_fd_sc_hd__nand3_4 _36822_ (.A(_14251_),
    .B(_14252_),
    .C(_14253_),
    .Y(_14254_));
 sky130_vsdinv _36823_ (.A(_13776_),
    .Y(_14255_));
 sky130_fd_sc_hd__a21o_2 _36824_ (.A1(_13769_),
    .A2(_13808_),
    .B1(_14255_),
    .X(_14256_));
 sky130_fd_sc_hd__and3_2 _36825_ (.A(_14250_),
    .B(_14254_),
    .C(_14256_),
    .X(_14257_));
 sky130_fd_sc_hd__a21oi_4 _36826_ (.A1(_14250_),
    .A2(_14254_),
    .B1(_14256_),
    .Y(_14258_));
 sky130_fd_sc_hd__o2bb2ai_4 _36827_ (.A1_N(_14183_),
    .A2_N(_14188_),
    .B1(_14257_),
    .B2(_14258_),
    .Y(_14259_));
 sky130_fd_sc_hd__nor2_4 _36828_ (.A(_14258_),
    .B(_14257_),
    .Y(_14260_));
 sky130_fd_sc_hd__nand3_4 _36829_ (.A(_14260_),
    .B(_14188_),
    .C(_14183_),
    .Y(_14261_));
 sky130_fd_sc_hd__a22oi_4 _36830_ (.A1(_14063_),
    .A2(_13953_),
    .B1(_14259_),
    .B2(_14261_),
    .Y(_14262_));
 sky130_fd_sc_hd__a21o_1 _36831_ (.A1(_14250_),
    .A2(_14254_),
    .B1(_14256_),
    .X(_14263_));
 sky130_fd_sc_hd__nand3_2 _36832_ (.A(_14250_),
    .B(_14254_),
    .C(_14256_),
    .Y(_14264_));
 sky130_fd_sc_hd__nand2_4 _36833_ (.A(_14263_),
    .B(_14264_),
    .Y(_14265_));
 sky130_fd_sc_hd__a21o_2 _36834_ (.A1(_14188_),
    .A2(_14183_),
    .B1(_14265_),
    .X(_14266_));
 sky130_fd_sc_hd__nand3_4 _36835_ (.A(_14188_),
    .B(_14265_),
    .C(_14183_),
    .Y(_14267_));
 sky130_fd_sc_hd__nand2_4 _36836_ (.A(_14063_),
    .B(_13953_),
    .Y(_14268_));
 sky130_fd_sc_hd__a21oi_4 _36837_ (.A1(_14266_),
    .A2(_14267_),
    .B1(_14268_),
    .Y(_14269_));
 sky130_vsdinv _36838_ (.A(_13978_),
    .Y(_14270_));
 sky130_vsdinv _36839_ (.A(_13974_),
    .Y(_14271_));
 sky130_fd_sc_hd__nor2_2 _36840_ (.A(_13979_),
    .B(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__a21oi_4 _36841_ (.A1(_13777_),
    .A2(_13778_),
    .B1(_13780_),
    .Y(_14273_));
 sky130_fd_sc_hd__nor2_2 _36842_ (.A(_13779_),
    .B(_14273_),
    .Y(_14274_));
 sky130_fd_sc_hd__nand3_4 _36843_ (.A(_14274_),
    .B(_13976_),
    .C(_13977_),
    .Y(_14275_));
 sky130_fd_sc_hd__o211ai_4 _36844_ (.A1(_13779_),
    .A2(_14273_),
    .B1(_13973_),
    .C1(_13970_),
    .Y(_14276_));
 sky130_fd_sc_hd__or2_1 _36845_ (.A(_13969_),
    .B(_13971_),
    .X(_14277_));
 sky130_fd_sc_hd__buf_2 _36846_ (.A(_14277_),
    .X(_14278_));
 sky130_fd_sc_hd__clkbuf_4 _36847_ (.A(_14278_),
    .X(_14279_));
 sky130_fd_sc_hd__a21o_2 _36848_ (.A1(_14275_),
    .A2(_14276_),
    .B1(_14279_),
    .X(_14280_));
 sky130_fd_sc_hd__nand3_4 _36849_ (.A(_14275_),
    .B(_14276_),
    .C(_14279_),
    .Y(_14281_));
 sky130_fd_sc_hd__a21oi_2 _36850_ (.A1(_13793_),
    .A2(_13797_),
    .B1(_13801_),
    .Y(_14282_));
 sky130_fd_sc_hd__o21ai_4 _36851_ (.A1(_13786_),
    .A2(_14282_),
    .B1(_13802_),
    .Y(_14283_));
 sky130_fd_sc_hd__a21oi_4 _36852_ (.A1(_14280_),
    .A2(_14281_),
    .B1(_14283_),
    .Y(_14284_));
 sky130_vsdinv _36853_ (.A(_14276_),
    .Y(_14285_));
 sky130_fd_sc_hd__buf_4 _36854_ (.A(_14277_),
    .X(_14286_));
 sky130_fd_sc_hd__nand2_1 _36855_ (.A(_14275_),
    .B(_14286_),
    .Y(_14287_));
 sky130_fd_sc_hd__o211a_1 _36856_ (.A1(_14285_),
    .A2(_14287_),
    .B1(_14280_),
    .C1(_14283_),
    .X(_14288_));
 sky130_fd_sc_hd__o22ai_4 _36857_ (.A1(_14270_),
    .A2(_14272_),
    .B1(_14284_),
    .B2(_14288_),
    .Y(_14289_));
 sky130_fd_sc_hd__a21oi_1 _36858_ (.A1(_13978_),
    .A2(_13979_),
    .B1(_14271_),
    .Y(_14290_));
 sky130_fd_sc_hd__a21o_1 _36859_ (.A1(_14280_),
    .A2(_14281_),
    .B1(_14283_),
    .X(_14291_));
 sky130_fd_sc_hd__nand3_4 _36860_ (.A(_14283_),
    .B(_14280_),
    .C(_14281_),
    .Y(_14292_));
 sky130_fd_sc_hd__nand3b_4 _36861_ (.A_N(_14290_),
    .B(_14291_),
    .C(_14292_),
    .Y(_14293_));
 sky130_fd_sc_hd__nand2_1 _36862_ (.A(_13983_),
    .B(_13989_),
    .Y(_14294_));
 sky130_fd_sc_hd__nand2_2 _36863_ (.A(_14294_),
    .B(_13987_),
    .Y(_14295_));
 sky130_fd_sc_hd__a21oi_4 _36864_ (.A1(_14289_),
    .A2(_14293_),
    .B1(_14295_),
    .Y(_14296_));
 sky130_fd_sc_hd__nor2_1 _36865_ (.A(_13982_),
    .B(_14000_),
    .Y(_14297_));
 sky130_fd_sc_hd__o211a_2 _36866_ (.A1(_14297_),
    .A2(_14001_),
    .B1(_14293_),
    .C1(_14289_),
    .X(_14298_));
 sky130_fd_sc_hd__o21ai_2 _36867_ (.A1(_14296_),
    .A2(_14298_),
    .B1(_13687_),
    .Y(_14299_));
 sky130_fd_sc_hd__nand2_1 _36868_ (.A(_13816_),
    .B(_13817_),
    .Y(_14300_));
 sky130_fd_sc_hd__nand2_2 _36869_ (.A(_14300_),
    .B(_13813_),
    .Y(_14301_));
 sky130_fd_sc_hd__a21o_1 _36870_ (.A1(_14289_),
    .A2(_14293_),
    .B1(_14295_),
    .X(_14302_));
 sky130_fd_sc_hd__buf_4 _36871_ (.A(_13678_),
    .X(_14303_));
 sky130_fd_sc_hd__nand3_2 _36872_ (.A(_14295_),
    .B(_14289_),
    .C(_14293_),
    .Y(_14304_));
 sky130_fd_sc_hd__nand3_2 _36873_ (.A(_14302_),
    .B(_14303_),
    .C(_14304_),
    .Y(_14305_));
 sky130_fd_sc_hd__nand3_4 _36874_ (.A(_14299_),
    .B(_14301_),
    .C(_14305_),
    .Y(_14306_));
 sky130_fd_sc_hd__o22ai_4 _36875_ (.A1(_13689_),
    .A2(_13675_),
    .B1(_14296_),
    .B2(_14298_),
    .Y(_14307_));
 sky130_fd_sc_hd__a22oi_2 _36876_ (.A1(_13524_),
    .A2(_13811_),
    .B1(_13805_),
    .B2(_13809_),
    .Y(_14308_));
 sky130_fd_sc_hd__o21ai_2 _36877_ (.A1(_13817_),
    .A2(_14308_),
    .B1(_13816_),
    .Y(_14309_));
 sky130_fd_sc_hd__buf_4 _36878_ (.A(_13677_),
    .X(_14310_));
 sky130_fd_sc_hd__nand3_2 _36879_ (.A(_14302_),
    .B(_14310_),
    .C(_14304_),
    .Y(_14311_));
 sky130_fd_sc_hd__nand3_4 _36880_ (.A(_14307_),
    .B(_14309_),
    .C(_14311_),
    .Y(_14312_));
 sky130_fd_sc_hd__nand2_1 _36881_ (.A(_14306_),
    .B(_14312_),
    .Y(_14313_));
 sky130_vsdinv _36882_ (.A(_14003_),
    .Y(_14314_));
 sky130_fd_sc_hd__a21o_1 _36883_ (.A1(_13687_),
    .A2(_13998_),
    .B1(_14314_),
    .X(_14315_));
 sky130_vsdinv _36884_ (.A(_14315_),
    .Y(_14316_));
 sky130_fd_sc_hd__nand2_1 _36885_ (.A(_14313_),
    .B(_14316_),
    .Y(_14317_));
 sky130_fd_sc_hd__nand3_4 _36886_ (.A(_14306_),
    .B(_14312_),
    .C(_14315_),
    .Y(_14318_));
 sky130_fd_sc_hd__and2_1 _36887_ (.A(_14317_),
    .B(_14318_),
    .X(_14319_));
 sky130_fd_sc_hd__o21ai_4 _36888_ (.A1(_14262_),
    .A2(_14269_),
    .B1(_14319_),
    .Y(_14320_));
 sky130_fd_sc_hd__nand3_4 _36889_ (.A(_14268_),
    .B(_14266_),
    .C(_14267_),
    .Y(_14321_));
 sky130_fd_sc_hd__o21ai_2 _36890_ (.A1(_13961_),
    .A2(_13949_),
    .B1(_13955_),
    .Y(_14322_));
 sky130_fd_sc_hd__nand3_4 _36891_ (.A(_14322_),
    .B(_14259_),
    .C(_14261_),
    .Y(_14323_));
 sky130_fd_sc_hd__nand2_4 _36892_ (.A(_14317_),
    .B(_14318_),
    .Y(_14324_));
 sky130_fd_sc_hd__nand3_4 _36893_ (.A(_14321_),
    .B(_14323_),
    .C(_14324_),
    .Y(_14325_));
 sky130_fd_sc_hd__nand3_4 _36894_ (.A(_14062_),
    .B(_14320_),
    .C(_14325_),
    .Y(_14326_));
 sky130_fd_sc_hd__nand2_2 _36895_ (.A(_14028_),
    .B(_13957_),
    .Y(_14327_));
 sky130_fd_sc_hd__a31oi_4 _36896_ (.A1(_14268_),
    .A2(_14267_),
    .A3(_14266_),
    .B1(_14324_),
    .Y(_14328_));
 sky130_fd_sc_hd__nand2_1 _36897_ (.A(_14328_),
    .B(_14323_),
    .Y(_14329_));
 sky130_fd_sc_hd__o21ai_2 _36898_ (.A1(_14262_),
    .A2(_14269_),
    .B1(_14324_),
    .Y(_14330_));
 sky130_fd_sc_hd__nand3_4 _36899_ (.A(_14327_),
    .B(_14329_),
    .C(_14330_),
    .Y(_14331_));
 sky130_fd_sc_hd__nand2_2 _36900_ (.A(_14021_),
    .B(_14017_),
    .Y(_14332_));
 sky130_fd_sc_hd__a21oi_4 _36901_ (.A1(_14332_),
    .A2(_14017_),
    .B1(_13740_),
    .Y(_14333_));
 sky130_fd_sc_hd__nand2_2 _36902_ (.A(_14017_),
    .B(_13740_),
    .Y(_14334_));
 sky130_fd_sc_hd__nor2_4 _36903_ (.A(_14334_),
    .B(_14018_),
    .Y(_14335_));
 sky130_fd_sc_hd__o2bb2ai_4 _36904_ (.A1_N(_14326_),
    .A2_N(_14331_),
    .B1(_14333_),
    .B2(_14335_),
    .Y(_14336_));
 sky130_fd_sc_hd__a21o_1 _36905_ (.A1(_14332_),
    .A2(_14017_),
    .B1(_13740_),
    .X(_14337_));
 sky130_fd_sc_hd__o21ai_2 _36906_ (.A1(_14018_),
    .A2(_14334_),
    .B1(_14337_),
    .Y(_14338_));
 sky130_fd_sc_hd__a31oi_4 _36907_ (.A1(_14062_),
    .A2(_14320_),
    .A3(_14325_),
    .B1(_14338_),
    .Y(_14339_));
 sky130_fd_sc_hd__nand2_2 _36908_ (.A(_14339_),
    .B(_14331_),
    .Y(_14340_));
 sky130_fd_sc_hd__o21ai_4 _36909_ (.A1(_14038_),
    .A2(_14026_),
    .B1(_14032_),
    .Y(_14341_));
 sky130_fd_sc_hd__a21oi_4 _36910_ (.A1(_14336_),
    .A2(_14340_),
    .B1(_14341_),
    .Y(_14342_));
 sky130_fd_sc_hd__a21oi_4 _36911_ (.A1(_14320_),
    .A2(_14325_),
    .B1(_14062_),
    .Y(_14343_));
 sky130_fd_sc_hd__nor2_2 _36912_ (.A(_14335_),
    .B(_14333_),
    .Y(_14344_));
 sky130_fd_sc_hd__nand2_1 _36913_ (.A(_14326_),
    .B(_14344_),
    .Y(_14345_));
 sky130_fd_sc_hd__o211a_1 _36914_ (.A1(_14343_),
    .A2(_14345_),
    .B1(_14336_),
    .C1(_14341_),
    .X(_14346_));
 sky130_fd_sc_hd__o21ai_1 _36915_ (.A1(_14342_),
    .A2(_14346_),
    .B1(_13744_),
    .Y(_14347_));
 sky130_fd_sc_hd__a21o_1 _36916_ (.A1(_14336_),
    .A2(_14340_),
    .B1(_14341_),
    .X(_14348_));
 sky130_vsdinv _36917_ (.A(_13744_),
    .Y(_14349_));
 sky130_fd_sc_hd__nand3_2 _36918_ (.A(_14341_),
    .B(_14336_),
    .C(_14340_),
    .Y(_14350_));
 sky130_fd_sc_hd__nand3_1 _36919_ (.A(_14348_),
    .B(_14349_),
    .C(_14350_),
    .Y(_14351_));
 sky130_fd_sc_hd__nand3b_2 _36920_ (.A_N(_14061_),
    .B(_14347_),
    .C(_14351_),
    .Y(_14352_));
 sky130_fd_sc_hd__clkbuf_8 _36921_ (.A(_13739_),
    .X(_14353_));
 sky130_fd_sc_hd__clkbuf_8 _36922_ (.A(_14353_),
    .X(_14354_));
 sky130_fd_sc_hd__buf_2 _36923_ (.A(_14354_),
    .X(_14355_));
 sky130_fd_sc_hd__clkbuf_4 _36924_ (.A(net412),
    .X(_14356_));
 sky130_fd_sc_hd__o22ai_1 _36925_ (.A1(_14356_),
    .A2(_13742_),
    .B1(_14342_),
    .B2(_14346_),
    .Y(_14357_));
 sky130_fd_sc_hd__nand3_1 _36926_ (.A(_14348_),
    .B(_13744_),
    .C(_14350_),
    .Y(_14358_));
 sky130_fd_sc_hd__nand3_2 _36927_ (.A(_14357_),
    .B(_14061_),
    .C(_14358_),
    .Y(_14359_));
 sky130_fd_sc_hd__and2_2 _36928_ (.A(_14352_),
    .B(_14359_),
    .X(_14360_));
 sky130_fd_sc_hd__nand2_2 _36929_ (.A(_14057_),
    .B(_14048_),
    .Y(_14361_));
 sky130_fd_sc_hd__xor2_4 _36930_ (.A(_14360_),
    .B(_14361_),
    .X(_02660_));
 sky130_fd_sc_hd__nand2_1 _36931_ (.A(_14081_),
    .B(_14082_),
    .Y(_14362_));
 sky130_fd_sc_hd__a21oi_2 _36932_ (.A1(_14083_),
    .A2(_14362_),
    .B1(_14092_),
    .Y(_14363_));
 sky130_fd_sc_hd__a22oi_4 _36933_ (.A1(_14363_),
    .A2(_14085_),
    .B1(_14093_),
    .B2(_14103_),
    .Y(_14364_));
 sky130_fd_sc_hd__nand2_2 _36934_ (.A(_19843_),
    .B(_06714_),
    .Y(_14365_));
 sky130_fd_sc_hd__nand2_4 _36935_ (.A(\pcpi_mul.rs2[29] ),
    .B(_06142_),
    .Y(_14366_));
 sky130_fd_sc_hd__nand2_4 _36936_ (.A(_19839_),
    .B(_06294_),
    .Y(_14367_));
 sky130_fd_sc_hd__nor2_8 _36937_ (.A(_14366_),
    .B(_14367_),
    .Y(_14368_));
 sky130_fd_sc_hd__and2_1 _36938_ (.A(_14366_),
    .B(_14367_),
    .X(_14369_));
 sky130_fd_sc_hd__nor2_2 _36939_ (.A(_14368_),
    .B(_14369_),
    .Y(_14370_));
 sky130_fd_sc_hd__nor2_2 _36940_ (.A(_14365_),
    .B(_14370_),
    .Y(_14371_));
 sky130_vsdinv _36941_ (.A(_14368_),
    .Y(_14372_));
 sky130_fd_sc_hd__nand2_4 _36942_ (.A(_14366_),
    .B(_14367_),
    .Y(_14373_));
 sky130_fd_sc_hd__and3_1 _36943_ (.A(_14372_),
    .B(_14365_),
    .C(_14373_),
    .X(_14374_));
 sky130_fd_sc_hd__nand3_2 _36944_ (.A(_11778_),
    .B(_11777_),
    .C(_05999_),
    .Y(_14375_));
 sky130_fd_sc_hd__nor2_2 _36945_ (.A(_10919_),
    .B(_14375_),
    .Y(_14376_));
 sky130_fd_sc_hd__a22oi_4 _36946_ (.A1(_10972_),
    .A2(_08530_),
    .B1(_06287_),
    .B2(_10973_),
    .Y(_14377_));
 sky130_fd_sc_hd__o22ai_4 _36947_ (.A1(net441),
    .A2(_07191_),
    .B1(_14376_),
    .B2(_14377_),
    .Y(_14378_));
 sky130_fd_sc_hd__nand2_1 _36948_ (.A(_19828_),
    .B(_07024_),
    .Y(_14379_));
 sky130_fd_sc_hd__nand3b_4 _36949_ (.A_N(_14379_),
    .B(_13139_),
    .C(net445),
    .Y(_14380_));
 sky130_fd_sc_hd__o21ai_2 _36950_ (.A1(_10919_),
    .A2(_13142_),
    .B1(_14379_),
    .Y(_14381_));
 sky130_fd_sc_hd__nand2_2 _36951_ (.A(_10573_),
    .B(_07185_),
    .Y(_14382_));
 sky130_vsdinv _36952_ (.A(_14382_),
    .Y(_14383_));
 sky130_fd_sc_hd__nand3_4 _36953_ (.A(_14380_),
    .B(_14381_),
    .C(_14383_),
    .Y(_14384_));
 sky130_fd_sc_hd__o22ai_4 _36954_ (.A1(net454),
    .A2(_14076_),
    .B1(_14083_),
    .B2(_14078_),
    .Y(_14385_));
 sky130_fd_sc_hd__a21oi_4 _36955_ (.A1(_14378_),
    .A2(_14384_),
    .B1(_14385_),
    .Y(_14386_));
 sky130_fd_sc_hd__o21ai_1 _36956_ (.A1(_20147_),
    .A2(_14375_),
    .B1(_14383_),
    .Y(_14387_));
 sky130_fd_sc_hd__o211a_4 _36957_ (.A1(_14377_),
    .A2(_14387_),
    .B1(_14385_),
    .C1(_14378_),
    .X(_14388_));
 sky130_fd_sc_hd__o22ai_4 _36958_ (.A1(_14371_),
    .A2(_14374_),
    .B1(_14386_),
    .B2(_14388_),
    .Y(_14389_));
 sky130_fd_sc_hd__a21o_2 _36959_ (.A1(_14378_),
    .A2(_14384_),
    .B1(_14385_),
    .X(_14390_));
 sky130_fd_sc_hd__nand3_4 _36960_ (.A(_14378_),
    .B(_14385_),
    .C(_14384_),
    .Y(_14391_));
 sky130_fd_sc_hd__inv_2 _36961_ (.A(_14365_),
    .Y(_14392_));
 sky130_fd_sc_hd__nand3_1 _36962_ (.A(_14372_),
    .B(_14392_),
    .C(_14373_),
    .Y(_14393_));
 sky130_fd_sc_hd__o21ai_1 _36963_ (.A1(_14368_),
    .A2(_14369_),
    .B1(_14365_),
    .Y(_14394_));
 sky130_fd_sc_hd__nand2_1 _36964_ (.A(_14393_),
    .B(_14394_),
    .Y(_14395_));
 sky130_fd_sc_hd__nand3_2 _36965_ (.A(_14390_),
    .B(_14391_),
    .C(_14395_),
    .Y(_14396_));
 sky130_fd_sc_hd__nand3_4 _36966_ (.A(_14364_),
    .B(_14389_),
    .C(_14396_),
    .Y(_14397_));
 sky130_fd_sc_hd__nor2_2 _36967_ (.A(_14392_),
    .B(_14370_),
    .Y(_14398_));
 sky130_fd_sc_hd__and3_1 _36968_ (.A(_14372_),
    .B(_14392_),
    .C(_14373_),
    .X(_14399_));
 sky130_fd_sc_hd__o22ai_4 _36969_ (.A1(_14398_),
    .A2(_14399_),
    .B1(_14386_),
    .B2(_14388_),
    .Y(_14400_));
 sky130_fd_sc_hd__o21ai_2 _36970_ (.A1(_14097_),
    .A2(_14087_),
    .B1(_14094_),
    .Y(_14401_));
 sky130_fd_sc_hd__nand3_1 _36971_ (.A(_14372_),
    .B(_14365_),
    .C(_14373_),
    .Y(_14402_));
 sky130_fd_sc_hd__o21ai_1 _36972_ (.A1(_14368_),
    .A2(_14369_),
    .B1(_14392_),
    .Y(_14403_));
 sky130_fd_sc_hd__nand2_2 _36973_ (.A(_14402_),
    .B(_14403_),
    .Y(_14404_));
 sky130_fd_sc_hd__nand3_4 _36974_ (.A(_14390_),
    .B(_14391_),
    .C(_14404_),
    .Y(_14405_));
 sky130_fd_sc_hd__nand3_2 _36975_ (.A(_14400_),
    .B(_14401_),
    .C(_14405_),
    .Y(_14406_));
 sky130_fd_sc_hd__buf_4 _36976_ (.A(_14406_),
    .X(_14407_));
 sky130_fd_sc_hd__nand2_1 _36977_ (.A(_14397_),
    .B(_14407_),
    .Y(_14408_));
 sky130_fd_sc_hd__and2_2 _36978_ (.A(_14112_),
    .B(_14108_),
    .X(_14409_));
 sky130_fd_sc_hd__nand2_2 _36979_ (.A(_09980_),
    .B(_07257_),
    .Y(_14410_));
 sky130_fd_sc_hd__a21o_1 _36980_ (.A1(_12818_),
    .A2(_07568_),
    .B1(_14410_),
    .X(_14411_));
 sky130_fd_sc_hd__nand2_1 _36981_ (.A(_19851_),
    .B(_20123_),
    .Y(_14412_));
 sky130_fd_sc_hd__a21o_1 _36982_ (.A1(_11366_),
    .A2(_10350_),
    .B1(_14412_),
    .X(_14413_));
 sky130_fd_sc_hd__nand2_2 _36983_ (.A(_08802_),
    .B(_07250_),
    .Y(_14414_));
 sky130_fd_sc_hd__nand3_4 _36984_ (.A(_14411_),
    .B(_14413_),
    .C(_14414_),
    .Y(_14415_));
 sky130_fd_sc_hd__nand3b_4 _36985_ (.A_N(_14410_),
    .B(_11010_),
    .C(_09443_),
    .Y(_14416_));
 sky130_vsdinv _36986_ (.A(_14414_),
    .Y(_14417_));
 sky130_fd_sc_hd__nand2_1 _36987_ (.A(_14410_),
    .B(_14412_),
    .Y(_14418_));
 sky130_fd_sc_hd__nand3_4 _36988_ (.A(_14416_),
    .B(_14417_),
    .C(_14418_),
    .Y(_14419_));
 sky130_fd_sc_hd__o21a_1 _36989_ (.A1(_14070_),
    .A2(_14071_),
    .B1(_14068_),
    .X(_14420_));
 sky130_fd_sc_hd__nor2_4 _36990_ (.A(_14069_),
    .B(_14420_),
    .Y(_14421_));
 sky130_fd_sc_hd__a21oi_4 _36991_ (.A1(_14415_),
    .A2(_14419_),
    .B1(_14421_),
    .Y(_14422_));
 sky130_fd_sc_hd__nor2_2 _36992_ (.A(_14409_),
    .B(_14422_),
    .Y(_14423_));
 sky130_fd_sc_hd__nand3_4 _36993_ (.A(_14421_),
    .B(_14415_),
    .C(_14419_),
    .Y(_14424_));
 sky130_fd_sc_hd__o2bb2ai_2 _36994_ (.A1_N(_14415_),
    .A2_N(_14419_),
    .B1(_14069_),
    .B2(_14420_),
    .Y(_14425_));
 sky130_fd_sc_hd__nand2_2 _36995_ (.A(_14112_),
    .B(_14108_),
    .Y(_14426_));
 sky130_fd_sc_hd__a21oi_4 _36996_ (.A1(_14425_),
    .A2(_14424_),
    .B1(_14426_),
    .Y(_14427_));
 sky130_fd_sc_hd__a21oi_4 _36997_ (.A1(_14423_),
    .A2(_14424_),
    .B1(_14427_),
    .Y(_14428_));
 sky130_fd_sc_hd__nand2_1 _36998_ (.A(_14408_),
    .B(_14428_),
    .Y(_14429_));
 sky130_fd_sc_hd__a21oi_2 _36999_ (.A1(_14090_),
    .A2(_14098_),
    .B1(_14067_),
    .Y(_14430_));
 sky130_fd_sc_hd__a21oi_2 _37000_ (.A1(_14099_),
    .A2(_14124_),
    .B1(_14430_),
    .Y(_14431_));
 sky130_fd_sc_hd__nor2_1 _37001_ (.A(_14068_),
    .B(_14069_),
    .Y(_14432_));
 sky130_fd_sc_hd__o211a_2 _37002_ (.A1(_14072_),
    .A2(_14432_),
    .B1(_14419_),
    .C1(_14415_),
    .X(_14433_));
 sky130_fd_sc_hd__nand2_2 _37003_ (.A(_14425_),
    .B(_14426_),
    .Y(_14434_));
 sky130_fd_sc_hd__o21ai_2 _37004_ (.A1(_14422_),
    .A2(_14433_),
    .B1(_14409_),
    .Y(_14435_));
 sky130_fd_sc_hd__o21ai_4 _37005_ (.A1(_14433_),
    .A2(_14434_),
    .B1(_14435_),
    .Y(_14436_));
 sky130_fd_sc_hd__nand3_2 _37006_ (.A(_14397_),
    .B(_14407_),
    .C(_14436_),
    .Y(_14437_));
 sky130_fd_sc_hd__nand3_4 _37007_ (.A(_14429_),
    .B(_14431_),
    .C(_14437_),
    .Y(_14438_));
 sky130_fd_sc_hd__nand2_2 _37008_ (.A(_14099_),
    .B(_14124_),
    .Y(_14439_));
 sky130_fd_sc_hd__nand2_2 _37009_ (.A(_14439_),
    .B(_14105_),
    .Y(_14440_));
 sky130_fd_sc_hd__nor2_2 _37010_ (.A(_14433_),
    .B(_14434_),
    .Y(_14441_));
 sky130_fd_sc_hd__o2bb2ai_4 _37011_ (.A1_N(_14407_),
    .A2_N(_14397_),
    .B1(_14427_),
    .B2(_14441_),
    .Y(_14442_));
 sky130_fd_sc_hd__nand3_4 _37012_ (.A(_14428_),
    .B(_14397_),
    .C(_14407_),
    .Y(_14443_));
 sky130_fd_sc_hd__nand3_4 _37013_ (.A(_14440_),
    .B(_14442_),
    .C(_14443_),
    .Y(_14444_));
 sky130_fd_sc_hd__o22ai_4 _37014_ (.A1(_12073_),
    .A2(_14139_),
    .B1(_14141_),
    .B2(_14138_),
    .Y(_14445_));
 sky130_fd_sc_hd__a22oi_4 _37015_ (.A1(_10917_),
    .A2(_08060_),
    .B1(_10926_),
    .B2(_10711_),
    .Y(_14446_));
 sky130_fd_sc_hd__nand3_4 _37016_ (.A(_10433_),
    .B(_07965_),
    .C(_07561_),
    .Y(_14447_));
 sky130_fd_sc_hd__nor2_4 _37017_ (.A(_10340_),
    .B(_14447_),
    .Y(_14448_));
 sky130_fd_sc_hd__nand2_4 _37018_ (.A(_19866_),
    .B(_08052_),
    .Y(_14449_));
 sky130_vsdinv _37019_ (.A(_14449_),
    .Y(_14450_));
 sky130_fd_sc_hd__o21ai_2 _37020_ (.A1(_14446_),
    .A2(_14448_),
    .B1(_14450_),
    .Y(_14451_));
 sky130_fd_sc_hd__a22o_2 _37021_ (.A1(_13902_),
    .A2(_10113_),
    .B1(_12447_),
    .B2(_10711_),
    .X(_14452_));
 sky130_fd_sc_hd__o211ai_4 _37022_ (.A1(_10340_),
    .A2(_14447_),
    .B1(_14449_),
    .C1(_14452_),
    .Y(_14453_));
 sky130_fd_sc_hd__nand3b_4 _37023_ (.A_N(_14445_),
    .B(_14451_),
    .C(_14453_),
    .Y(_14454_));
 sky130_fd_sc_hd__o21ai_2 _37024_ (.A1(_14446_),
    .A2(_14448_),
    .B1(_14449_),
    .Y(_14455_));
 sky130_fd_sc_hd__o211ai_2 _37025_ (.A1(_10824_),
    .A2(_14447_),
    .B1(_14450_),
    .C1(_14452_),
    .Y(_14456_));
 sky130_fd_sc_hd__nand3_4 _37026_ (.A(_14455_),
    .B(_14456_),
    .C(_14445_),
    .Y(_14457_));
 sky130_fd_sc_hd__nand2_2 _37027_ (.A(_10628_),
    .B(_20104_),
    .Y(_14458_));
 sky130_fd_sc_hd__nand2_2 _37028_ (.A(_10944_),
    .B(_20101_),
    .Y(_14459_));
 sky130_fd_sc_hd__nor2_2 _37029_ (.A(_14458_),
    .B(_14459_),
    .Y(_14460_));
 sky130_fd_sc_hd__and2_1 _37030_ (.A(_14458_),
    .B(_14459_),
    .X(_14461_));
 sky130_fd_sc_hd__nand2_1 _37031_ (.A(_11869_),
    .B(_12103_),
    .Y(_14462_));
 sky130_vsdinv _37032_ (.A(_14462_),
    .Y(_14463_));
 sky130_fd_sc_hd__o21ai_1 _37033_ (.A1(_14460_),
    .A2(_14461_),
    .B1(_14463_),
    .Y(_14464_));
 sky130_fd_sc_hd__nand2_1 _37034_ (.A(_14458_),
    .B(_14459_),
    .Y(_14465_));
 sky130_fd_sc_hd__nand3b_1 _37035_ (.A_N(_14460_),
    .B(_14462_),
    .C(_14465_),
    .Y(_14466_));
 sky130_fd_sc_hd__nand2_2 _37036_ (.A(_14464_),
    .B(_14466_),
    .Y(_14467_));
 sky130_fd_sc_hd__a21o_2 _37037_ (.A1(_14454_),
    .A2(_14457_),
    .B1(_14467_),
    .X(_14468_));
 sky130_fd_sc_hd__nand3_4 _37038_ (.A(_14467_),
    .B(_14454_),
    .C(_14457_),
    .Y(_14469_));
 sky130_fd_sc_hd__and2_1 _37039_ (.A(_13875_),
    .B(_13872_),
    .X(_14470_));
 sky130_fd_sc_hd__o21ai_4 _37040_ (.A1(_14117_),
    .A2(_14470_),
    .B1(_14119_),
    .Y(_14471_));
 sky130_fd_sc_hd__a21o_2 _37041_ (.A1(_14468_),
    .A2(_14469_),
    .B1(_14471_),
    .X(_14472_));
 sky130_fd_sc_hd__nand3_4 _37042_ (.A(_14471_),
    .B(_14468_),
    .C(_14469_),
    .Y(_14473_));
 sky130_fd_sc_hd__nand2_4 _37043_ (.A(_14170_),
    .B(_14149_),
    .Y(_14474_));
 sky130_fd_sc_hd__a21oi_4 _37044_ (.A1(_14472_),
    .A2(_14473_),
    .B1(_14474_),
    .Y(_14475_));
 sky130_vsdinv _37045_ (.A(_14457_),
    .Y(_14476_));
 sky130_fd_sc_hd__nand2_1 _37046_ (.A(_14467_),
    .B(_14454_),
    .Y(_14477_));
 sky130_fd_sc_hd__o211a_2 _37047_ (.A1(_14476_),
    .A2(_14477_),
    .B1(_14468_),
    .C1(_14471_),
    .X(_14478_));
 sky130_fd_sc_hd__nand2_2 _37048_ (.A(_14472_),
    .B(_14474_),
    .Y(_14479_));
 sky130_fd_sc_hd__nor2_4 _37049_ (.A(_14478_),
    .B(_14479_),
    .Y(_14480_));
 sky130_fd_sc_hd__o2bb2ai_4 _37050_ (.A1_N(_14438_),
    .A2_N(_14444_),
    .B1(_14475_),
    .B2(_14480_),
    .Y(_14481_));
 sky130_vsdinv _37051_ (.A(_14149_),
    .Y(_14482_));
 sky130_fd_sc_hd__a21oi_4 _37052_ (.A1(_14468_),
    .A2(_14469_),
    .B1(_14471_),
    .Y(_14483_));
 sky130_fd_sc_hd__o22ai_4 _37053_ (.A1(_14482_),
    .A2(_14164_),
    .B1(_14483_),
    .B2(_14478_),
    .Y(_14484_));
 sky130_vsdinv _37054_ (.A(_14474_),
    .Y(_14485_));
 sky130_fd_sc_hd__nand3_2 _37055_ (.A(_14472_),
    .B(_14485_),
    .C(_14473_),
    .Y(_14486_));
 sky130_fd_sc_hd__nand2_4 _37056_ (.A(_14484_),
    .B(_14486_),
    .Y(_14487_));
 sky130_fd_sc_hd__nand3_4 _37057_ (.A(_14438_),
    .B(_14444_),
    .C(_14487_),
    .Y(_14488_));
 sky130_vsdinv _37058_ (.A(_14134_),
    .Y(_14489_));
 sky130_fd_sc_hd__nand2_1 _37059_ (.A(_14131_),
    .B(_14133_),
    .Y(_14490_));
 sky130_fd_sc_hd__o2bb2ai_4 _37060_ (.A1_N(_14181_),
    .A2_N(_14130_),
    .B1(_14489_),
    .B2(_14490_),
    .Y(_14491_));
 sky130_fd_sc_hd__a21oi_4 _37061_ (.A1(_14481_),
    .A2(_14488_),
    .B1(_14491_),
    .Y(_14492_));
 sky130_fd_sc_hd__and3_1 _37062_ (.A(_14440_),
    .B(_14442_),
    .C(_14443_),
    .X(_14493_));
 sky130_fd_sc_hd__nand2_1 _37063_ (.A(_14438_),
    .B(_14487_),
    .Y(_14494_));
 sky130_fd_sc_hd__o211a_1 _37064_ (.A1(_14493_),
    .A2(_14494_),
    .B1(_14491_),
    .C1(_14481_),
    .X(_14495_));
 sky130_vsdinv _37065_ (.A(_14205_),
    .Y(_14496_));
 sky130_fd_sc_hd__and3_1 _37066_ (.A(_14194_),
    .B(_14199_),
    .C(_14197_),
    .X(_14497_));
 sky130_fd_sc_hd__nor2_2 _37067_ (.A(_14206_),
    .B(_14497_),
    .Y(_14498_));
 sky130_fd_sc_hd__nand2_2 _37068_ (.A(_07754_),
    .B(_09037_),
    .Y(_14499_));
 sky130_fd_sc_hd__nand3_2 _37069_ (.A(_14499_),
    .B(_19888_),
    .C(_13456_),
    .Y(_14500_));
 sky130_fd_sc_hd__a21o_1 _37070_ (.A1(_19888_),
    .A2(_11927_),
    .B1(_14499_),
    .X(_14501_));
 sky130_fd_sc_hd__o211ai_4 _37071_ (.A1(net443),
    .A2(_12307_),
    .B1(_14500_),
    .C1(_14501_),
    .Y(_14502_));
 sky130_fd_sc_hd__nand3b_4 _37072_ (.A_N(_14499_),
    .B(_12576_),
    .C(_11210_),
    .Y(_14503_));
 sky130_fd_sc_hd__nor2_2 _37073_ (.A(_06528_),
    .B(_10265_),
    .Y(_14504_));
 sky130_fd_sc_hd__a22o_1 _37074_ (.A1(_19881_),
    .A2(_09038_),
    .B1(_07090_),
    .B2(_20090_),
    .X(_14505_));
 sky130_fd_sc_hd__nand3_4 _37075_ (.A(_14503_),
    .B(_14504_),
    .C(_14505_),
    .Y(_14506_));
 sky130_fd_sc_hd__nor2_2 _37076_ (.A(_14158_),
    .B(_14156_),
    .Y(_14507_));
 sky130_fd_sc_hd__o2bb2ai_4 _37077_ (.A1_N(_14502_),
    .A2_N(_14506_),
    .B1(_14155_),
    .B2(_14507_),
    .Y(_14508_));
 sky130_fd_sc_hd__o21bai_4 _37078_ (.A1(_14157_),
    .A2(_14155_),
    .B1_N(_14156_),
    .Y(_14509_));
 sky130_fd_sc_hd__nand3_4 _37079_ (.A(_14509_),
    .B(_14502_),
    .C(_14506_),
    .Y(_14510_));
 sky130_fd_sc_hd__nor2_2 _37080_ (.A(_14193_),
    .B(_14190_),
    .Y(_14511_));
 sky130_fd_sc_hd__nor2_2 _37081_ (.A(_14192_),
    .B(_14511_),
    .Y(_14512_));
 sky130_vsdinv _37082_ (.A(_14512_),
    .Y(_14513_));
 sky130_fd_sc_hd__a21oi_2 _37083_ (.A1(_14508_),
    .A2(_14510_),
    .B1(_14513_),
    .Y(_14514_));
 sky130_fd_sc_hd__o211a_1 _37084_ (.A1(_14192_),
    .A2(_14511_),
    .B1(_14510_),
    .C1(_14508_),
    .X(_14515_));
 sky130_fd_sc_hd__o22ai_4 _37085_ (.A1(_14496_),
    .A2(_14498_),
    .B1(_14514_),
    .B2(_14515_),
    .Y(_14516_));
 sky130_fd_sc_hd__a21bo_2 _37086_ (.A1(_14206_),
    .A2(_14205_),
    .B1_N(_14200_),
    .X(_14517_));
 sky130_fd_sc_hd__nor2_2 _37087_ (.A(_14195_),
    .B(_14192_),
    .Y(_14518_));
 sky130_fd_sc_hd__a21oi_4 _37088_ (.A1(_14502_),
    .A2(_14506_),
    .B1(_14509_),
    .Y(_14519_));
 sky130_fd_sc_hd__nor2_1 _37089_ (.A(_14157_),
    .B(_14155_),
    .Y(_14520_));
 sky130_fd_sc_hd__o211a_1 _37090_ (.A1(_14156_),
    .A2(_14520_),
    .B1(_14506_),
    .C1(_14502_),
    .X(_14521_));
 sky130_fd_sc_hd__o22ai_4 _37091_ (.A1(_14190_),
    .A2(_14518_),
    .B1(_14519_),
    .B2(_14521_),
    .Y(_14522_));
 sky130_fd_sc_hd__nand3_4 _37092_ (.A(_14508_),
    .B(_14513_),
    .C(_14510_),
    .Y(_14523_));
 sky130_fd_sc_hd__nand3_4 _37093_ (.A(_14517_),
    .B(_14522_),
    .C(_14523_),
    .Y(_14524_));
 sky130_fd_sc_hd__nand2_4 _37094_ (.A(_07102_),
    .B(\pcpi_mul.rs1[28] ),
    .Y(_14525_));
 sky130_fd_sc_hd__nand3b_2 _37095_ (.A_N(_14525_),
    .B(_10693_),
    .C(_10761_),
    .Y(_14526_));
 sky130_fd_sc_hd__nor2_4 _37096_ (.A(_13271_),
    .B(_10766_),
    .Y(_14527_));
 sky130_fd_sc_hd__nand2_4 _37097_ (.A(_06607_),
    .B(_20077_),
    .Y(_14528_));
 sky130_fd_sc_hd__nand2_4 _37098_ (.A(_14525_),
    .B(_14528_),
    .Y(_14529_));
 sky130_fd_sc_hd__nand3_4 _37099_ (.A(_14526_),
    .B(_14527_),
    .C(_14529_),
    .Y(_14530_));
 sky130_fd_sc_hd__nand3_2 _37100_ (.A(_14528_),
    .B(_10692_),
    .C(_09896_),
    .Y(_14531_));
 sky130_fd_sc_hd__nand3_2 _37101_ (.A(_14525_),
    .B(_06208_),
    .C(_20078_),
    .Y(_14532_));
 sky130_fd_sc_hd__o211ai_4 _37102_ (.A1(_13271_),
    .A2(_10766_),
    .B1(_14531_),
    .C1(_14532_),
    .Y(_14533_));
 sky130_fd_sc_hd__nand2_4 _37103_ (.A(_14530_),
    .B(_14533_),
    .Y(_14534_));
 sky130_fd_sc_hd__a21oi_4 _37104_ (.A1(_14221_),
    .A2(_14220_),
    .B1(_14217_),
    .Y(_14535_));
 sky130_fd_sc_hd__nand2_1 _37105_ (.A(_14534_),
    .B(_14535_),
    .Y(_14536_));
 sky130_fd_sc_hd__a21o_1 _37106_ (.A1(_14221_),
    .A2(_14220_),
    .B1(_14217_),
    .X(_14537_));
 sky130_fd_sc_hd__nand3_4 _37107_ (.A(_14537_),
    .B(_14533_),
    .C(_14530_),
    .Y(_14538_));
 sky130_fd_sc_hd__nand2_4 _37108_ (.A(_06630_),
    .B(\pcpi_mul.rs1[31] ),
    .Y(_14539_));
 sky130_fd_sc_hd__nand2_8 _37109_ (.A(net504),
    .B(_06534_),
    .Y(_14540_));
 sky130_fd_sc_hd__nor2_8 _37110_ (.A(_14539_),
    .B(_14540_),
    .Y(_14541_));
 sky130_fd_sc_hd__and2_1 _37111_ (.A(_14539_),
    .B(_14540_),
    .X(_14542_));
 sky130_fd_sc_hd__o21ai_2 _37112_ (.A1(_14541_),
    .A2(_14542_),
    .B1(_14235_),
    .Y(_14543_));
 sky130_fd_sc_hd__nand2_1 _37113_ (.A(_14539_),
    .B(_14540_),
    .Y(_14544_));
 sky130_fd_sc_hd__nand3b_4 _37114_ (.A_N(_14541_),
    .B(_14234_),
    .C(_14544_),
    .Y(_14545_));
 sky130_fd_sc_hd__nand2_1 _37115_ (.A(_14543_),
    .B(_14545_),
    .Y(_14546_));
 sky130_fd_sc_hd__a21o_1 _37116_ (.A1(_14536_),
    .A2(_14538_),
    .B1(_14546_),
    .X(_14547_));
 sky130_fd_sc_hd__a22oi_4 _37117_ (.A1(_14543_),
    .A2(_14545_),
    .B1(_14534_),
    .B2(_14535_),
    .Y(_14548_));
 sky130_fd_sc_hd__nand2_1 _37118_ (.A(_14548_),
    .B(_14538_),
    .Y(_14549_));
 sky130_fd_sc_hd__nand2_2 _37119_ (.A(_14547_),
    .B(_14549_),
    .Y(_14550_));
 sky130_fd_sc_hd__a21boi_4 _37120_ (.A1(_14516_),
    .A2(_14524_),
    .B1_N(_14550_),
    .Y(_14551_));
 sky130_fd_sc_hd__a21oi_4 _37121_ (.A1(_14522_),
    .A2(_14523_),
    .B1(_14517_),
    .Y(_14552_));
 sky130_fd_sc_hd__o211a_4 _37122_ (.A1(_14497_),
    .A2(_14212_),
    .B1(_14523_),
    .C1(_14522_),
    .X(_14553_));
 sky130_fd_sc_hd__nor3_4 _37123_ (.A(_14550_),
    .B(_14552_),
    .C(_14553_),
    .Y(_14554_));
 sky130_fd_sc_hd__nand2_4 _37124_ (.A(_14175_),
    .B(_14171_),
    .Y(_14555_));
 sky130_fd_sc_hd__o21bai_4 _37125_ (.A1(_14551_),
    .A2(_14554_),
    .B1_N(_14555_),
    .Y(_14556_));
 sky130_fd_sc_hd__a21oi_2 _37126_ (.A1(_14536_),
    .A2(_14538_),
    .B1(_14546_),
    .Y(_14557_));
 sky130_vsdinv _37127_ (.A(_14549_),
    .Y(_14558_));
 sky130_fd_sc_hd__o22ai_4 _37128_ (.A1(_14557_),
    .A2(_14558_),
    .B1(_14552_),
    .B2(_14553_),
    .Y(_14559_));
 sky130_fd_sc_hd__nand3b_4 _37129_ (.A_N(_14550_),
    .B(_14516_),
    .C(_14524_),
    .Y(_14560_));
 sky130_fd_sc_hd__nand3_4 _37130_ (.A(_14559_),
    .B(_14555_),
    .C(_14560_),
    .Y(_14561_));
 sky130_fd_sc_hd__a21oi_4 _37131_ (.A1(_14211_),
    .A2(_14213_),
    .B1(_14210_),
    .Y(_14562_));
 sky130_fd_sc_hd__nor2_2 _37132_ (.A(_14247_),
    .B(_14248_),
    .Y(_14563_));
 sky130_fd_sc_hd__o21ai_4 _37133_ (.A1(_14562_),
    .A2(_14563_),
    .B1(_14214_),
    .Y(_14564_));
 sky130_fd_sc_hd__a21oi_4 _37134_ (.A1(_14556_),
    .A2(_14561_),
    .B1(_14564_),
    .Y(_14565_));
 sky130_vsdinv _37135_ (.A(_14564_),
    .Y(_14566_));
 sky130_fd_sc_hd__a21oi_4 _37136_ (.A1(_14559_),
    .A2(_14560_),
    .B1(_14555_),
    .Y(_14567_));
 sky130_fd_sc_hd__o211a_2 _37137_ (.A1(_14174_),
    .A2(_14180_),
    .B1(_14560_),
    .C1(_14559_),
    .X(_14568_));
 sky130_fd_sc_hd__nor3_4 _37138_ (.A(_14566_),
    .B(_14567_),
    .C(_14568_),
    .Y(_14569_));
 sky130_fd_sc_hd__nor2_4 _37139_ (.A(_14565_),
    .B(_14569_),
    .Y(_14570_));
 sky130_fd_sc_hd__o21ai_2 _37140_ (.A1(_14492_),
    .A2(_14495_),
    .B1(_14570_),
    .Y(_14571_));
 sky130_fd_sc_hd__a21boi_4 _37141_ (.A1(_14260_),
    .A2(_14188_),
    .B1_N(_14183_),
    .Y(_14572_));
 sky130_fd_sc_hd__a21oi_1 _37142_ (.A1(_14438_),
    .A2(_14444_),
    .B1(_14487_),
    .Y(_14573_));
 sky130_fd_sc_hd__and3_1 _37143_ (.A(_14438_),
    .B(_14444_),
    .C(_14487_),
    .X(_14574_));
 sky130_fd_sc_hd__o21bai_2 _37144_ (.A1(_14573_),
    .A2(_14574_),
    .B1_N(_14491_),
    .Y(_14575_));
 sky130_fd_sc_hd__nand3_4 _37145_ (.A(_14481_),
    .B(_14491_),
    .C(_14488_),
    .Y(_14576_));
 sky130_fd_sc_hd__o21bai_2 _37146_ (.A1(_14567_),
    .A2(_14568_),
    .B1_N(_14564_),
    .Y(_14577_));
 sky130_fd_sc_hd__nand3_2 _37147_ (.A(_14556_),
    .B(_14564_),
    .C(_14561_),
    .Y(_14578_));
 sky130_fd_sc_hd__nand2_4 _37148_ (.A(_14577_),
    .B(_14578_),
    .Y(_14579_));
 sky130_fd_sc_hd__nand3_2 _37149_ (.A(_14575_),
    .B(_14576_),
    .C(_14579_),
    .Y(_14580_));
 sky130_fd_sc_hd__nand3_4 _37150_ (.A(_14571_),
    .B(_14572_),
    .C(_14580_),
    .Y(_14581_));
 sky130_fd_sc_hd__o22ai_4 _37151_ (.A1(_14569_),
    .A2(_14565_),
    .B1(_14492_),
    .B2(_14495_),
    .Y(_14582_));
 sky130_fd_sc_hd__a21oi_4 _37152_ (.A1(_14177_),
    .A2(_14182_),
    .B1(_14066_),
    .Y(_14583_));
 sky130_fd_sc_hd__o21ai_4 _37153_ (.A1(_14265_),
    .A2(_14583_),
    .B1(_14183_),
    .Y(_14584_));
 sky130_fd_sc_hd__nand3_4 _37154_ (.A(_14570_),
    .B(_14575_),
    .C(_14576_),
    .Y(_14585_));
 sky130_fd_sc_hd__nand3_4 _37155_ (.A(_14582_),
    .B(_14584_),
    .C(_14585_),
    .Y(_14586_));
 sky130_fd_sc_hd__nand2_1 _37156_ (.A(_14581_),
    .B(_14586_),
    .Y(_14587_));
 sky130_fd_sc_hd__a21oi_4 _37157_ (.A1(_14230_),
    .A2(_14231_),
    .B1(_14234_),
    .Y(_14588_));
 sky130_fd_sc_hd__nor2_2 _37158_ (.A(_14232_),
    .B(_14588_),
    .Y(_14589_));
 sky130_fd_sc_hd__nand3_4 _37159_ (.A(_14589_),
    .B(_13976_),
    .C(_13977_),
    .Y(_14590_));
 sky130_fd_sc_hd__o211ai_4 _37160_ (.A1(_14232_),
    .A2(_14588_),
    .B1(_13973_),
    .C1(_13970_),
    .Y(_14591_));
 sky130_fd_sc_hd__a21oi_1 _37161_ (.A1(_14590_),
    .A2(_14591_),
    .B1(_14279_),
    .Y(_14592_));
 sky130_fd_sc_hd__and3_1 _37162_ (.A(_14590_),
    .B(_14591_),
    .C(_14286_),
    .X(_14593_));
 sky130_fd_sc_hd__a21oi_2 _37163_ (.A1(_14239_),
    .A2(_14237_),
    .B1(_14228_),
    .Y(_14594_));
 sky130_fd_sc_hd__o21ai_2 _37164_ (.A1(_14592_),
    .A2(_14593_),
    .B1(_14594_),
    .Y(_14595_));
 sky130_vsdinv _37165_ (.A(_14222_),
    .Y(_14596_));
 sky130_fd_sc_hd__nand2_1 _37166_ (.A(_14224_),
    .B(_14219_),
    .Y(_14597_));
 sky130_fd_sc_hd__o22ai_4 _37167_ (.A1(_14596_),
    .A2(_14597_),
    .B1(_14243_),
    .B2(_14225_),
    .Y(_14598_));
 sky130_fd_sc_hd__nand3_4 _37168_ (.A(_14590_),
    .B(_14591_),
    .C(_14279_),
    .Y(_14599_));
 sky130_fd_sc_hd__a21o_1 _37169_ (.A1(_14590_),
    .A2(_14591_),
    .B1(_14279_),
    .X(_14600_));
 sky130_fd_sc_hd__nand3_4 _37170_ (.A(_14598_),
    .B(_14599_),
    .C(_14600_),
    .Y(_14601_));
 sky130_fd_sc_hd__nand2_2 _37171_ (.A(_14287_),
    .B(_14276_),
    .Y(_14602_));
 sky130_fd_sc_hd__a21o_1 _37172_ (.A1(_14595_),
    .A2(_14601_),
    .B1(_14602_),
    .X(_14603_));
 sky130_fd_sc_hd__o21ai_1 _37173_ (.A1(_14290_),
    .A2(_14284_),
    .B1(_14292_),
    .Y(_14604_));
 sky130_fd_sc_hd__nand3_1 _37174_ (.A(_14595_),
    .B(_14601_),
    .C(_14602_),
    .Y(_14605_));
 sky130_fd_sc_hd__nand3_1 _37175_ (.A(_14603_),
    .B(_14604_),
    .C(_14605_),
    .Y(_14606_));
 sky130_fd_sc_hd__clkbuf_4 _37176_ (.A(_14606_),
    .X(_14607_));
 sky130_fd_sc_hd__a21oi_2 _37177_ (.A1(_14595_),
    .A2(_14601_),
    .B1(_14602_),
    .Y(_14608_));
 sky130_vsdinv _37178_ (.A(_14287_),
    .Y(_14609_));
 sky130_fd_sc_hd__o211a_1 _37179_ (.A1(_14285_),
    .A2(_14609_),
    .B1(_14601_),
    .C1(_14595_),
    .X(_14610_));
 sky130_fd_sc_hd__o21bai_4 _37180_ (.A1(_14608_),
    .A2(_14610_),
    .B1_N(_14604_),
    .Y(_14611_));
 sky130_fd_sc_hd__o2bb2ai_4 _37181_ (.A1_N(_14607_),
    .A2_N(_14611_),
    .B1(_13689_),
    .B2(_13675_),
    .Y(_14612_));
 sky130_fd_sc_hd__nand3_4 _37182_ (.A(_14611_),
    .B(_14009_),
    .C(_14607_),
    .Y(_14613_));
 sky130_fd_sc_hd__and2_1 _37183_ (.A(_13808_),
    .B(_13769_),
    .X(_14614_));
 sky130_fd_sc_hd__nor2_2 _37184_ (.A(_14255_),
    .B(_14614_),
    .Y(_14615_));
 sky130_fd_sc_hd__a21oi_2 _37185_ (.A1(_14252_),
    .A2(_14253_),
    .B1(_14251_),
    .Y(_14616_));
 sky130_fd_sc_hd__o21ai_4 _37186_ (.A1(_14615_),
    .A2(_14616_),
    .B1(_14254_),
    .Y(_14617_));
 sky130_fd_sc_hd__a21oi_4 _37187_ (.A1(_14612_),
    .A2(_14613_),
    .B1(_14617_),
    .Y(_14618_));
 sky130_vsdinv _37188_ (.A(_14607_),
    .Y(_14619_));
 sky130_fd_sc_hd__nand2_1 _37189_ (.A(_14611_),
    .B(_13687_),
    .Y(_14620_));
 sky130_fd_sc_hd__o211a_1 _37190_ (.A1(_14619_),
    .A2(_14620_),
    .B1(_14612_),
    .C1(_14617_),
    .X(_14621_));
 sky130_fd_sc_hd__a21oi_4 _37191_ (.A1(_14302_),
    .A2(_14014_),
    .B1(_14298_),
    .Y(_14622_));
 sky130_fd_sc_hd__o21ai_2 _37192_ (.A1(_14618_),
    .A2(_14621_),
    .B1(_14622_),
    .Y(_14623_));
 sky130_fd_sc_hd__a21oi_2 _37193_ (.A1(_14611_),
    .A2(_14607_),
    .B1(_14014_),
    .Y(_14624_));
 sky130_fd_sc_hd__and3_1 _37194_ (.A(_14611_),
    .B(_14310_),
    .C(_14606_),
    .X(_14625_));
 sky130_fd_sc_hd__o21bai_4 _37195_ (.A1(_14624_),
    .A2(_14625_),
    .B1_N(_14617_),
    .Y(_14626_));
 sky130_fd_sc_hd__nand3_4 _37196_ (.A(_14617_),
    .B(_14612_),
    .C(_14613_),
    .Y(_14627_));
 sky130_fd_sc_hd__nand3b_4 _37197_ (.A_N(_14622_),
    .B(_14626_),
    .C(_14627_),
    .Y(_14628_));
 sky130_fd_sc_hd__nand2_4 _37198_ (.A(_14623_),
    .B(_14628_),
    .Y(_14629_));
 sky130_fd_sc_hd__nand2_1 _37199_ (.A(_14319_),
    .B(_14321_),
    .Y(_14630_));
 sky130_fd_sc_hd__a22oi_4 _37200_ (.A1(_14587_),
    .A2(_14629_),
    .B1(_14630_),
    .B2(_14323_),
    .Y(_14631_));
 sky130_fd_sc_hd__a21boi_4 _37201_ (.A1(_14626_),
    .A2(_14627_),
    .B1_N(_14622_),
    .Y(_14632_));
 sky130_fd_sc_hd__nor3_4 _37202_ (.A(_14622_),
    .B(_14618_),
    .C(_14621_),
    .Y(_14633_));
 sky130_fd_sc_hd__nor2_2 _37203_ (.A(_14632_),
    .B(_14633_),
    .Y(_14634_));
 sky130_fd_sc_hd__nand3_4 _37204_ (.A(_14634_),
    .B(_14586_),
    .C(_14581_),
    .Y(_14635_));
 sky130_fd_sc_hd__nand2_2 _37205_ (.A(_14631_),
    .B(_14635_),
    .Y(_14636_));
 sky130_fd_sc_hd__o2bb2ai_4 _37206_ (.A1_N(_14586_),
    .A2_N(_14581_),
    .B1(_14632_),
    .B2(_14633_),
    .Y(_14637_));
 sky130_fd_sc_hd__nand2_1 _37207_ (.A(_14637_),
    .B(_14635_),
    .Y(_14638_));
 sky130_fd_sc_hd__nor2_2 _37208_ (.A(_14269_),
    .B(_14328_),
    .Y(_14639_));
 sky130_fd_sc_hd__nand2_4 _37209_ (.A(_14638_),
    .B(_14639_),
    .Y(_14640_));
 sky130_vsdinv _37210_ (.A(_13739_),
    .Y(_14641_));
 sky130_fd_sc_hd__and3_2 _37211_ (.A(_14318_),
    .B(_14641_),
    .C(_14312_),
    .X(_14642_));
 sky130_fd_sc_hd__and2_4 _37212_ (.A(_14318_),
    .B(_14312_),
    .X(_14643_));
 sky130_fd_sc_hd__nor2_8 _37213_ (.A(_14641_),
    .B(_14643_),
    .Y(_14644_));
 sky130_fd_sc_hd__nor2_8 _37214_ (.A(_14642_),
    .B(_14644_),
    .Y(_14645_));
 sky130_vsdinv _37215_ (.A(_14645_),
    .Y(_14646_));
 sky130_fd_sc_hd__nand3_4 _37216_ (.A(_14636_),
    .B(_14640_),
    .C(_14646_),
    .Y(_14647_));
 sky130_fd_sc_hd__o21ai_2 _37217_ (.A1(_14324_),
    .A2(_14262_),
    .B1(_14323_),
    .Y(_14648_));
 sky130_fd_sc_hd__a21oi_4 _37218_ (.A1(_14637_),
    .A2(_14635_),
    .B1(_14648_),
    .Y(_14649_));
 sky130_fd_sc_hd__o211a_1 _37219_ (.A1(_14269_),
    .A2(_14328_),
    .B1(_14635_),
    .C1(_14637_),
    .X(_14650_));
 sky130_fd_sc_hd__o21ai_2 _37220_ (.A1(_14649_),
    .A2(_14650_),
    .B1(_14645_),
    .Y(_14651_));
 sky130_fd_sc_hd__o211ai_4 _37221_ (.A1(_14343_),
    .A2(_14339_),
    .B1(_14647_),
    .C1(_14651_),
    .Y(_14652_));
 sky130_fd_sc_hd__o22ai_4 _37222_ (.A1(_14644_),
    .A2(_14642_),
    .B1(_14649_),
    .B2(_14650_),
    .Y(_14653_));
 sky130_fd_sc_hd__a21oi_2 _37223_ (.A1(_14326_),
    .A2(_14344_),
    .B1(_14343_),
    .Y(_14654_));
 sky130_fd_sc_hd__nand3_2 _37224_ (.A(_14636_),
    .B(_14640_),
    .C(_14645_),
    .Y(_14655_));
 sky130_fd_sc_hd__nand3_4 _37225_ (.A(_14653_),
    .B(_14654_),
    .C(_14655_),
    .Y(_14656_));
 sky130_fd_sc_hd__a21oi_1 _37226_ (.A1(_14652_),
    .A2(_14656_),
    .B1(_14333_),
    .Y(_14657_));
 sky130_fd_sc_hd__and3_1 _37227_ (.A(_14652_),
    .B(_14656_),
    .C(_14333_),
    .X(_14658_));
 sky130_fd_sc_hd__a21oi_1 _37228_ (.A1(_14348_),
    .A2(_13744_),
    .B1(_14346_),
    .Y(_14659_));
 sky130_fd_sc_hd__o21ai_2 _37229_ (.A1(_14657_),
    .A2(_14658_),
    .B1(_14659_),
    .Y(_14660_));
 sky130_fd_sc_hd__o21ai_2 _37230_ (.A1(_14349_),
    .A2(_14342_),
    .B1(_14350_),
    .Y(_14661_));
 sky130_fd_sc_hd__nand2_1 _37231_ (.A(_14652_),
    .B(_14656_),
    .Y(_14662_));
 sky130_fd_sc_hd__nand2_1 _37232_ (.A(_14662_),
    .B(_14337_),
    .Y(_14663_));
 sky130_fd_sc_hd__nand3_2 _37233_ (.A(_14652_),
    .B(_14656_),
    .C(_14333_),
    .Y(_14664_));
 sky130_fd_sc_hd__nand3_4 _37234_ (.A(_14661_),
    .B(_14663_),
    .C(_14664_),
    .Y(_14665_));
 sky130_fd_sc_hd__and2_1 _37235_ (.A(_14660_),
    .B(_14665_),
    .X(_14666_));
 sky130_fd_sc_hd__nand2_2 _37236_ (.A(_14352_),
    .B(_14359_),
    .Y(_14667_));
 sky130_fd_sc_hd__nand2_1 _37237_ (.A(_14359_),
    .B(_14048_),
    .Y(_14668_));
 sky130_fd_sc_hd__nand2_1 _37238_ (.A(_14668_),
    .B(_14352_),
    .Y(_14669_));
 sky130_fd_sc_hd__o31ai_2 _37239_ (.A1(_14049_),
    .A2(_14667_),
    .A3(_14056_),
    .B1(_14669_),
    .Y(_14670_));
 sky130_fd_sc_hd__or2_1 _37240_ (.A(_14666_),
    .B(_14670_),
    .X(_14671_));
 sky130_fd_sc_hd__nand2_1 _37241_ (.A(_14670_),
    .B(_14666_),
    .Y(_14672_));
 sky130_fd_sc_hd__and2_4 _37242_ (.A(_14671_),
    .B(_14672_),
    .X(_02661_));
 sky130_fd_sc_hd__a22oi_4 _37243_ (.A1(_14635_),
    .A2(_14631_),
    .B1(_14640_),
    .B2(_14646_),
    .Y(_14673_));
 sky130_fd_sc_hd__nand2_4 _37244_ (.A(_14628_),
    .B(_14627_),
    .Y(_14674_));
 sky130_fd_sc_hd__nand2_1 _37245_ (.A(_14674_),
    .B(_13739_),
    .Y(_14675_));
 sky130_vsdinv _37246_ (.A(_14675_),
    .Y(_14676_));
 sky130_fd_sc_hd__nor2_8 _37247_ (.A(_14353_),
    .B(_14674_),
    .Y(_14677_));
 sky130_fd_sc_hd__o21ai_2 _37248_ (.A1(_14579_),
    .A2(_14492_),
    .B1(_14576_),
    .Y(_14678_));
 sky130_fd_sc_hd__nand2_2 _37249_ (.A(_14494_),
    .B(_14444_),
    .Y(_14679_));
 sky130_fd_sc_hd__a21oi_4 _37250_ (.A1(_14390_),
    .A2(_14404_),
    .B1(_14388_),
    .Y(_14680_));
 sky130_fd_sc_hd__nand2_2 _37251_ (.A(_09320_),
    .B(_07543_),
    .Y(_14681_));
 sky130_fd_sc_hd__a22oi_4 _37252_ (.A1(_10411_),
    .A2(_06718_),
    .B1(_10412_),
    .B2(_20130_),
    .Y(_14682_));
 sky130_fd_sc_hd__nand2_2 _37253_ (.A(_09996_),
    .B(_06437_),
    .Y(_14683_));
 sky130_fd_sc_hd__nand2_2 _37254_ (.A(_10000_),
    .B(_08002_),
    .Y(_14684_));
 sky130_fd_sc_hd__nor2_2 _37255_ (.A(_14683_),
    .B(_14684_),
    .Y(_14685_));
 sky130_fd_sc_hd__nor2_2 _37256_ (.A(_14682_),
    .B(_14685_),
    .Y(_14686_));
 sky130_fd_sc_hd__nor2_2 _37257_ (.A(_14681_),
    .B(_14686_),
    .Y(_14687_));
 sky130_fd_sc_hd__and2_1 _37258_ (.A(_14686_),
    .B(_14681_),
    .X(_14688_));
 sky130_fd_sc_hd__nand3_4 _37259_ (.A(_18693_),
    .B(_11777_),
    .C(_05986_),
    .Y(_14689_));
 sky130_fd_sc_hd__nor2_4 _37260_ (.A(_08008_),
    .B(_14689_),
    .Y(_14690_));
 sky130_fd_sc_hd__a22oi_4 _37261_ (.A1(_19829_),
    .A2(net466),
    .B1(_06307_),
    .B2(_12487_),
    .Y(_14691_));
 sky130_fd_sc_hd__o22ai_4 _37262_ (.A1(net441),
    .A2(_07510_),
    .B1(_14690_),
    .B2(_14691_),
    .Y(_14692_));
 sky130_fd_sc_hd__nand2_2 _37263_ (.A(_10575_),
    .B(_07502_),
    .Y(_14693_));
 sky130_fd_sc_hd__nand3b_4 _37264_ (.A_N(_14693_),
    .B(_13139_),
    .C(_06307_),
    .Y(_14694_));
 sky130_fd_sc_hd__o21ai_4 _37265_ (.A1(_08008_),
    .A2(_10968_),
    .B1(_14693_),
    .Y(_14695_));
 sky130_fd_sc_hd__nand2_2 _37266_ (.A(_10573_),
    .B(_06442_),
    .Y(_14696_));
 sky130_vsdinv _37267_ (.A(_14696_),
    .Y(_14697_));
 sky130_fd_sc_hd__nand3_4 _37268_ (.A(_14694_),
    .B(_14695_),
    .C(_14697_),
    .Y(_14698_));
 sky130_fd_sc_hd__o21ai_4 _37269_ (.A1(_14382_),
    .A2(_14377_),
    .B1(_14380_),
    .Y(_14699_));
 sky130_fd_sc_hd__a21oi_4 _37270_ (.A1(_14692_),
    .A2(_14698_),
    .B1(_14699_),
    .Y(_14700_));
 sky130_fd_sc_hd__o21ai_1 _37271_ (.A1(_20143_),
    .A2(_14689_),
    .B1(_14697_),
    .Y(_14701_));
 sky130_fd_sc_hd__o211a_1 _37272_ (.A1(_14691_),
    .A2(_14701_),
    .B1(_14699_),
    .C1(_14692_),
    .X(_14702_));
 sky130_fd_sc_hd__o22ai_4 _37273_ (.A1(_14687_),
    .A2(_14688_),
    .B1(_14700_),
    .B2(_14702_),
    .Y(_14703_));
 sky130_fd_sc_hd__a21o_1 _37274_ (.A1(_14692_),
    .A2(_14698_),
    .B1(_14699_),
    .X(_14704_));
 sky130_fd_sc_hd__nand3_4 _37275_ (.A(_14692_),
    .B(_14699_),
    .C(_14698_),
    .Y(_14705_));
 sky130_vsdinv _37276_ (.A(_14681_),
    .Y(_14706_));
 sky130_fd_sc_hd__nand2_1 _37277_ (.A(_14686_),
    .B(_14706_),
    .Y(_14707_));
 sky130_fd_sc_hd__o21ai_2 _37278_ (.A1(_14682_),
    .A2(_14685_),
    .B1(_14681_),
    .Y(_14708_));
 sky130_fd_sc_hd__nand2_4 _37279_ (.A(_14707_),
    .B(_14708_),
    .Y(_14709_));
 sky130_fd_sc_hd__nand3_2 _37280_ (.A(_14704_),
    .B(_14705_),
    .C(_14709_),
    .Y(_14710_));
 sky130_fd_sc_hd__nand3_4 _37281_ (.A(_14680_),
    .B(_14703_),
    .C(_14710_),
    .Y(_14711_));
 sky130_fd_sc_hd__o21ai_2 _37282_ (.A1(_14700_),
    .A2(_14702_),
    .B1(_14709_),
    .Y(_14712_));
 sky130_fd_sc_hd__o21ai_2 _37283_ (.A1(_14395_),
    .A2(_14386_),
    .B1(_14391_),
    .Y(_14713_));
 sky130_fd_sc_hd__nand3b_2 _37284_ (.A_N(_14709_),
    .B(_14704_),
    .C(_14705_),
    .Y(_14714_));
 sky130_fd_sc_hd__nand3_4 _37285_ (.A(_14712_),
    .B(_14713_),
    .C(_14714_),
    .Y(_14715_));
 sky130_fd_sc_hd__nand2_4 _37286_ (.A(_19847_),
    .B(_06979_),
    .Y(_14716_));
 sky130_fd_sc_hd__nand3_2 _37287_ (.A(_14716_),
    .B(_11363_),
    .C(_20119_),
    .Y(_14717_));
 sky130_fd_sc_hd__a21o_1 _37288_ (.A1(_11371_),
    .A2(_20119_),
    .B1(_14716_),
    .X(_14718_));
 sky130_fd_sc_hd__o211ai_4 _37289_ (.A1(_08615_),
    .A2(_12073_),
    .B1(_14717_),
    .C1(_14718_),
    .Y(_14719_));
 sky130_fd_sc_hd__nand3b_4 _37290_ (.A_N(_14716_),
    .B(_11371_),
    .C(_11061_),
    .Y(_14720_));
 sky130_fd_sc_hd__nor2_2 _37291_ (.A(net464),
    .B(_11057_),
    .Y(_14721_));
 sky130_fd_sc_hd__a22o_1 _37292_ (.A1(_19848_),
    .A2(_20123_),
    .B1(_11010_),
    .B2(_12059_),
    .X(_14722_));
 sky130_fd_sc_hd__nand3_4 _37293_ (.A(_14720_),
    .B(_14721_),
    .C(_14722_),
    .Y(_14723_));
 sky130_fd_sc_hd__nand2_2 _37294_ (.A(_14719_),
    .B(_14723_),
    .Y(_14724_));
 sky130_fd_sc_hd__a21oi_4 _37295_ (.A1(_14392_),
    .A2(_14373_),
    .B1(_14368_),
    .Y(_14725_));
 sky130_fd_sc_hd__nand2_1 _37296_ (.A(_14724_),
    .B(_14725_),
    .Y(_14726_));
 sky130_fd_sc_hd__a21o_2 _37297_ (.A1(_14392_),
    .A2(_14373_),
    .B1(_14368_),
    .X(_14727_));
 sky130_fd_sc_hd__nand3_4 _37298_ (.A(_14727_),
    .B(_14719_),
    .C(_14723_),
    .Y(_14728_));
 sky130_fd_sc_hd__and2_1 _37299_ (.A(_14419_),
    .B(_14416_),
    .X(_14729_));
 sky130_fd_sc_hd__a21boi_4 _37300_ (.A1(_14726_),
    .A2(_14728_),
    .B1_N(_14729_),
    .Y(_14730_));
 sky130_fd_sc_hd__a22oi_4 _37301_ (.A1(_14416_),
    .A2(_14419_),
    .B1(_14724_),
    .B2(_14725_),
    .Y(_14731_));
 sky130_fd_sc_hd__and2_1 _37302_ (.A(_14731_),
    .B(_14728_),
    .X(_14732_));
 sky130_fd_sc_hd__o2bb2ai_2 _37303_ (.A1_N(_14711_),
    .A2_N(_14715_),
    .B1(_14730_),
    .B2(_14732_),
    .Y(_14733_));
 sky130_fd_sc_hd__a21oi_4 _37304_ (.A1(_14400_),
    .A2(_14405_),
    .B1(_14401_),
    .Y(_14734_));
 sky130_fd_sc_hd__a21oi_4 _37305_ (.A1(_14407_),
    .A2(_14436_),
    .B1(_14734_),
    .Y(_14735_));
 sky130_fd_sc_hd__a21oi_4 _37306_ (.A1(_14728_),
    .A2(_14731_),
    .B1(_14730_),
    .Y(_14736_));
 sky130_fd_sc_hd__nand3_2 _37307_ (.A(_14736_),
    .B(_14711_),
    .C(_14715_),
    .Y(_14737_));
 sky130_fd_sc_hd__nand3_4 _37308_ (.A(_14733_),
    .B(_14735_),
    .C(_14737_),
    .Y(_14738_));
 sky130_fd_sc_hd__nand2_1 _37309_ (.A(_14711_),
    .B(_14715_),
    .Y(_14739_));
 sky130_fd_sc_hd__nand2_2 _37310_ (.A(_14739_),
    .B(_14736_),
    .Y(_14740_));
 sky130_fd_sc_hd__nand2_1 _37311_ (.A(_14406_),
    .B(_14436_),
    .Y(_14741_));
 sky130_fd_sc_hd__nand2_4 _37312_ (.A(_14741_),
    .B(_14397_),
    .Y(_14742_));
 sky130_fd_sc_hd__o211ai_4 _37313_ (.A1(_14730_),
    .A2(_14732_),
    .B1(_14715_),
    .C1(_14711_),
    .Y(_14743_));
 sky130_fd_sc_hd__nand3_4 _37314_ (.A(_14740_),
    .B(_14742_),
    .C(_14743_),
    .Y(_14744_));
 sky130_fd_sc_hd__a22oi_4 _37315_ (.A1(_19859_),
    .A2(_20111_),
    .B1(_10918_),
    .B2(_20108_),
    .Y(_14745_));
 sky130_fd_sc_hd__nand3_4 _37316_ (.A(_10440_),
    .B(_19863_),
    .C(_11487_),
    .Y(_14746_));
 sky130_fd_sc_hd__nor2_4 _37317_ (.A(_11734_),
    .B(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__nand2_4 _37318_ (.A(_19866_),
    .B(_09926_),
    .Y(_14748_));
 sky130_vsdinv _37319_ (.A(_14748_),
    .Y(_14749_));
 sky130_fd_sc_hd__o21ai_2 _37320_ (.A1(_14745_),
    .A2(_14747_),
    .B1(_14749_),
    .Y(_14750_));
 sky130_fd_sc_hd__a21oi_4 _37321_ (.A1(_14452_),
    .A2(_14450_),
    .B1(_14448_),
    .Y(_14751_));
 sky130_fd_sc_hd__a22o_1 _37322_ (.A1(_19859_),
    .A2(_10711_),
    .B1(_10918_),
    .B2(_10343_),
    .X(_14752_));
 sky130_fd_sc_hd__o211ai_2 _37323_ (.A1(_12093_),
    .A2(_14746_),
    .B1(_14748_),
    .C1(_14752_),
    .Y(_14753_));
 sky130_fd_sc_hd__nand3_4 _37324_ (.A(_14750_),
    .B(_14751_),
    .C(_14753_),
    .Y(_14754_));
 sky130_fd_sc_hd__o21ai_2 _37325_ (.A1(_14745_),
    .A2(_14747_),
    .B1(_14748_),
    .Y(_14755_));
 sky130_fd_sc_hd__o22ai_4 _37326_ (.A1(_10824_),
    .A2(_14447_),
    .B1(_14449_),
    .B2(_14446_),
    .Y(_14756_));
 sky130_fd_sc_hd__o211ai_2 _37327_ (.A1(_12093_),
    .A2(_14746_),
    .B1(_14749_),
    .C1(_14752_),
    .Y(_14757_));
 sky130_fd_sc_hd__nand3_4 _37328_ (.A(_14755_),
    .B(_14756_),
    .C(_14757_),
    .Y(_14758_));
 sky130_fd_sc_hd__nand2_2 _37329_ (.A(_19870_),
    .B(_08881_),
    .Y(_14759_));
 sky130_fd_sc_hd__nand2_2 _37330_ (.A(_07902_),
    .B(_12103_),
    .Y(_14760_));
 sky130_fd_sc_hd__nor2_1 _37331_ (.A(_14759_),
    .B(_14760_),
    .Y(_14761_));
 sky130_fd_sc_hd__and2_1 _37332_ (.A(_14759_),
    .B(_14760_),
    .X(_14762_));
 sky130_fd_sc_hd__nand2_2 _37333_ (.A(_11869_),
    .B(_10814_),
    .Y(_14763_));
 sky130_fd_sc_hd__o21bai_1 _37334_ (.A1(_14761_),
    .A2(_14762_),
    .B1_N(_14763_),
    .Y(_14764_));
 sky130_fd_sc_hd__nand2_1 _37335_ (.A(_14759_),
    .B(_14760_),
    .Y(_14765_));
 sky130_fd_sc_hd__nand3b_2 _37336_ (.A_N(_14761_),
    .B(_14763_),
    .C(_14765_),
    .Y(_14766_));
 sky130_fd_sc_hd__nand2_2 _37337_ (.A(_14764_),
    .B(_14766_),
    .Y(_14767_));
 sky130_fd_sc_hd__a21o_2 _37338_ (.A1(_14754_),
    .A2(_14758_),
    .B1(_14767_),
    .X(_14768_));
 sky130_fd_sc_hd__nand3_4 _37339_ (.A(_14767_),
    .B(_14754_),
    .C(_14758_),
    .Y(_14769_));
 sky130_fd_sc_hd__a21oi_4 _37340_ (.A1(_14409_),
    .A2(_14424_),
    .B1(_14422_),
    .Y(_14770_));
 sky130_fd_sc_hd__a21o_1 _37341_ (.A1(_14768_),
    .A2(_14769_),
    .B1(_14770_),
    .X(_14771_));
 sky130_fd_sc_hd__nand3_4 _37342_ (.A(_14770_),
    .B(_14768_),
    .C(_14769_),
    .Y(_14772_));
 sky130_fd_sc_hd__nand2_2 _37343_ (.A(_14477_),
    .B(_14457_),
    .Y(_14773_));
 sky130_fd_sc_hd__a21oi_4 _37344_ (.A1(_14771_),
    .A2(_14772_),
    .B1(_14773_),
    .Y(_14774_));
 sky130_vsdinv _37345_ (.A(_14773_),
    .Y(_14775_));
 sky130_fd_sc_hd__nand2_2 _37346_ (.A(_14771_),
    .B(_14772_),
    .Y(_14776_));
 sky130_fd_sc_hd__nor2_4 _37347_ (.A(_14775_),
    .B(_14776_),
    .Y(_14777_));
 sky130_fd_sc_hd__o2bb2ai_2 _37348_ (.A1_N(_14738_),
    .A2_N(_14744_),
    .B1(_14774_),
    .B2(_14777_),
    .Y(_14778_));
 sky130_fd_sc_hd__a21oi_4 _37349_ (.A1(_14768_),
    .A2(_14769_),
    .B1(_14770_),
    .Y(_14779_));
 sky130_fd_sc_hd__nor2_2 _37350_ (.A(_14775_),
    .B(_14779_),
    .Y(_14780_));
 sky130_fd_sc_hd__a21oi_4 _37351_ (.A1(_14772_),
    .A2(_14780_),
    .B1(_14774_),
    .Y(_14781_));
 sky130_fd_sc_hd__nand3_4 _37352_ (.A(_14781_),
    .B(_14744_),
    .C(_14738_),
    .Y(_14782_));
 sky130_fd_sc_hd__nand3_4 _37353_ (.A(_14679_),
    .B(_14778_),
    .C(_14782_),
    .Y(_14783_));
 sky130_fd_sc_hd__nor2_2 _37354_ (.A(_14773_),
    .B(_14776_),
    .Y(_14784_));
 sky130_fd_sc_hd__and2_1 _37355_ (.A(_14776_),
    .B(_14773_),
    .X(_14785_));
 sky130_fd_sc_hd__o2bb2ai_4 _37356_ (.A1_N(_14738_),
    .A2_N(_14744_),
    .B1(_14784_),
    .B2(_14785_),
    .Y(_14786_));
 sky130_fd_sc_hd__a32oi_4 _37357_ (.A1(_14407_),
    .A2(_14397_),
    .A3(_14428_),
    .B1(_14439_),
    .B2(_14105_),
    .Y(_14787_));
 sky130_fd_sc_hd__a22oi_4 _37358_ (.A1(_14787_),
    .A2(_14442_),
    .B1(_14438_),
    .B2(_14487_),
    .Y(_14788_));
 sky130_fd_sc_hd__o211ai_4 _37359_ (.A1(_14774_),
    .A2(_14777_),
    .B1(_14744_),
    .C1(_14738_),
    .Y(_14789_));
 sky130_fd_sc_hd__nand3_4 _37360_ (.A(_14786_),
    .B(_14788_),
    .C(_14789_),
    .Y(_14790_));
 sky130_fd_sc_hd__nand2_1 _37361_ (.A(_14783_),
    .B(_14790_),
    .Y(_14791_));
 sky130_fd_sc_hd__nand2_2 _37362_ (.A(_11058_),
    .B(_10256_),
    .Y(_14792_));
 sky130_fd_sc_hd__a21o_1 _37363_ (.A1(_06360_),
    .A2(_10760_),
    .B1(_14792_),
    .X(_14793_));
 sky130_fd_sc_hd__nand2_2 _37364_ (.A(_06546_),
    .B(_11173_),
    .Y(_14794_));
 sky130_fd_sc_hd__a21o_1 _37365_ (.A1(_06369_),
    .A2(_10768_),
    .B1(_14794_),
    .X(_14795_));
 sky130_fd_sc_hd__o211ai_4 _37366_ (.A1(_13271_),
    .A2(_11177_),
    .B1(_14793_),
    .C1(_14795_),
    .Y(_14796_));
 sky130_fd_sc_hd__nand3_2 _37367_ (.A(_06369_),
    .B(_06360_),
    .C(_10768_),
    .Y(_14797_));
 sky130_fd_sc_hd__nand2_2 _37368_ (.A(_14792_),
    .B(_14794_),
    .Y(_14798_));
 sky130_fd_sc_hd__o2111ai_4 _37369_ (.A1(_10772_),
    .A2(_14797_),
    .B1(net455),
    .C1(_20070_),
    .D1(_14798_),
    .Y(_14799_));
 sky130_fd_sc_hd__nand2_1 _37370_ (.A(_14796_),
    .B(_14799_),
    .Y(_14800_));
 sky130_fd_sc_hd__nor2_2 _37371_ (.A(_14525_),
    .B(_14528_),
    .Y(_14801_));
 sky130_fd_sc_hd__a21oi_4 _37372_ (.A1(_14527_),
    .A2(_14529_),
    .B1(_14801_),
    .Y(_14802_));
 sky130_fd_sc_hd__nand2_2 _37373_ (.A(_14800_),
    .B(_14802_),
    .Y(_14803_));
 sky130_fd_sc_hd__a31o_2 _37374_ (.A1(_14529_),
    .A2(net455),
    .A3(_11607_),
    .B1(_14801_),
    .X(_14804_));
 sky130_fd_sc_hd__nand3_4 _37375_ (.A(_14804_),
    .B(_14799_),
    .C(_14796_),
    .Y(_14805_));
 sky130_fd_sc_hd__clkbuf_4 _37376_ (.A(\pcpi_mul.rs1[32] ),
    .X(_14806_));
 sky130_fd_sc_hd__o21a_1 _37377_ (.A1(_06344_),
    .A2(_06909_),
    .B1(_14806_),
    .X(_14807_));
 sky130_fd_sc_hd__nand3_4 _37378_ (.A(_14806_),
    .B(_06344_),
    .C(_05657_),
    .Y(_14808_));
 sky130_fd_sc_hd__nand2_4 _37379_ (.A(_14807_),
    .B(_14808_),
    .Y(_14809_));
 sky130_fd_sc_hd__nand2_2 _37380_ (.A(_14809_),
    .B(_14234_),
    .Y(_14810_));
 sky130_fd_sc_hd__o21a_2 _37381_ (.A1(_05633_),
    .A2(_14809_),
    .B1(_14810_),
    .X(_14811_));
 sky130_fd_sc_hd__clkbuf_4 _37382_ (.A(_14811_),
    .X(_14812_));
 sky130_fd_sc_hd__a21oi_4 _37383_ (.A1(_14803_),
    .A2(_14805_),
    .B1(_14812_),
    .Y(_14813_));
 sky130_fd_sc_hd__nand3_2 _37384_ (.A(_14803_),
    .B(_14805_),
    .C(_14812_),
    .Y(_14814_));
 sky130_vsdinv _37385_ (.A(_14814_),
    .Y(_14815_));
 sky130_fd_sc_hd__nand2_2 _37386_ (.A(_07289_),
    .B(_09025_),
    .Y(_14816_));
 sky130_fd_sc_hd__a21o_1 _37387_ (.A1(_06638_),
    .A2(_11934_),
    .B1(_14816_),
    .X(_14817_));
 sky130_fd_sc_hd__nand2_1 _37388_ (.A(_12576_),
    .B(_09899_),
    .Y(_14818_));
 sky130_fd_sc_hd__a21o_1 _37389_ (.A1(_11463_),
    .A2(_09902_),
    .B1(_14818_),
    .X(_14819_));
 sky130_fd_sc_hd__nand2_2 _37390_ (.A(_06641_),
    .B(_09896_),
    .Y(_14820_));
 sky130_fd_sc_hd__nand3_4 _37391_ (.A(_14817_),
    .B(_14819_),
    .C(_14820_),
    .Y(_14821_));
 sky130_fd_sc_hd__nand3b_4 _37392_ (.A_N(_14816_),
    .B(_11455_),
    .C(_11934_),
    .Y(_14822_));
 sky130_vsdinv _37393_ (.A(_14820_),
    .Y(_14823_));
 sky130_fd_sc_hd__nand2_1 _37394_ (.A(_14816_),
    .B(_14818_),
    .Y(_14824_));
 sky130_fd_sc_hd__nand3_4 _37395_ (.A(_14822_),
    .B(_14823_),
    .C(_14824_),
    .Y(_14825_));
 sky130_fd_sc_hd__a21o_2 _37396_ (.A1(_14463_),
    .A2(_14465_),
    .B1(_14460_),
    .X(_14826_));
 sky130_fd_sc_hd__a21oi_4 _37397_ (.A1(_14821_),
    .A2(_14825_),
    .B1(_14826_),
    .Y(_14827_));
 sky130_fd_sc_hd__a21oi_1 _37398_ (.A1(_14458_),
    .A2(_14459_),
    .B1(_14462_),
    .Y(_14828_));
 sky130_fd_sc_hd__o211a_1 _37399_ (.A1(_14460_),
    .A2(_14828_),
    .B1(_14825_),
    .C1(_14821_),
    .X(_14829_));
 sky130_fd_sc_hd__and2_2 _37400_ (.A(_14506_),
    .B(_14503_),
    .X(_14830_));
 sky130_fd_sc_hd__o21ai_4 _37401_ (.A1(_14827_),
    .A2(_14829_),
    .B1(_14830_),
    .Y(_14831_));
 sky130_fd_sc_hd__a21o_1 _37402_ (.A1(_14821_),
    .A2(_14825_),
    .B1(_14826_),
    .X(_14832_));
 sky130_fd_sc_hd__nand3_4 _37403_ (.A(_14826_),
    .B(_14821_),
    .C(_14825_),
    .Y(_14833_));
 sky130_fd_sc_hd__nand2_2 _37404_ (.A(_14506_),
    .B(_14503_),
    .Y(_14834_));
 sky130_fd_sc_hd__nand3_4 _37405_ (.A(_14832_),
    .B(_14833_),
    .C(_14834_),
    .Y(_14835_));
 sky130_fd_sc_hd__o21ai_4 _37406_ (.A1(_14512_),
    .A2(_14519_),
    .B1(_14510_),
    .Y(_14836_));
 sky130_fd_sc_hd__a21oi_4 _37407_ (.A1(_14831_),
    .A2(_14835_),
    .B1(_14836_),
    .Y(_14837_));
 sky130_fd_sc_hd__nand2_1 _37408_ (.A(_14832_),
    .B(_14834_),
    .Y(_14838_));
 sky130_fd_sc_hd__o211a_2 _37409_ (.A1(_14829_),
    .A2(_14838_),
    .B1(_14836_),
    .C1(_14831_),
    .X(_14839_));
 sky130_fd_sc_hd__o22ai_4 _37410_ (.A1(_14813_),
    .A2(_14815_),
    .B1(_14837_),
    .B2(_14839_),
    .Y(_14840_));
 sky130_fd_sc_hd__a21oi_4 _37411_ (.A1(_14796_),
    .A2(_14799_),
    .B1(_14804_),
    .Y(_14841_));
 sky130_fd_sc_hd__nor2_2 _37412_ (.A(_14802_),
    .B(_14800_),
    .Y(_14842_));
 sky130_fd_sc_hd__o21ai_4 _37413_ (.A1(_05633_),
    .A2(_14809_),
    .B1(_14810_),
    .Y(_14843_));
 sky130_fd_sc_hd__buf_4 _37414_ (.A(_14843_),
    .X(_14844_));
 sky130_fd_sc_hd__o21ai_1 _37415_ (.A1(_14841_),
    .A2(_14842_),
    .B1(_14844_),
    .Y(_14845_));
 sky130_fd_sc_hd__nand2_2 _37416_ (.A(_14845_),
    .B(_14814_),
    .Y(_14846_));
 sky130_fd_sc_hd__a21o_1 _37417_ (.A1(_14831_),
    .A2(_14835_),
    .B1(_14836_),
    .X(_14847_));
 sky130_fd_sc_hd__nand3_2 _37418_ (.A(_14831_),
    .B(_14835_),
    .C(_14836_),
    .Y(_14848_));
 sky130_fd_sc_hd__nand3b_4 _37419_ (.A_N(_14846_),
    .B(_14847_),
    .C(_14848_),
    .Y(_14849_));
 sky130_fd_sc_hd__nand2_2 _37420_ (.A(_14479_),
    .B(_14473_),
    .Y(_14850_));
 sky130_fd_sc_hd__a21oi_4 _37421_ (.A1(_14840_),
    .A2(_14849_),
    .B1(_14850_),
    .Y(_14851_));
 sky130_fd_sc_hd__nor2_1 _37422_ (.A(_14485_),
    .B(_14483_),
    .Y(_14852_));
 sky130_fd_sc_hd__o211a_2 _37423_ (.A1(_14478_),
    .A2(_14852_),
    .B1(_14849_),
    .C1(_14840_),
    .X(_14853_));
 sky130_fd_sc_hd__nor2_2 _37424_ (.A(_14550_),
    .B(_14552_),
    .Y(_14854_));
 sky130_fd_sc_hd__nor2_4 _37425_ (.A(_14553_),
    .B(_14854_),
    .Y(_14855_));
 sky130_fd_sc_hd__o21ai_4 _37426_ (.A1(_14851_),
    .A2(_14853_),
    .B1(_14855_),
    .Y(_14856_));
 sky130_vsdinv _37427_ (.A(_14855_),
    .Y(_14857_));
 sky130_fd_sc_hd__nor2_2 _37428_ (.A(_14474_),
    .B(_14478_),
    .Y(_14858_));
 sky130_fd_sc_hd__o2bb2ai_4 _37429_ (.A1_N(_14849_),
    .A2_N(_14840_),
    .B1(_14483_),
    .B2(_14858_),
    .Y(_14859_));
 sky130_fd_sc_hd__nand3_4 _37430_ (.A(_14850_),
    .B(_14849_),
    .C(_14840_),
    .Y(_14860_));
 sky130_fd_sc_hd__nand3_4 _37431_ (.A(_14857_),
    .B(_14859_),
    .C(_14860_),
    .Y(_14861_));
 sky130_fd_sc_hd__nand2_1 _37432_ (.A(_14856_),
    .B(_14861_),
    .Y(_14862_));
 sky130_fd_sc_hd__nand2_2 _37433_ (.A(_14791_),
    .B(_14862_),
    .Y(_14863_));
 sky130_fd_sc_hd__a21oi_1 _37434_ (.A1(_14859_),
    .A2(_14860_),
    .B1(_14857_),
    .Y(_14864_));
 sky130_fd_sc_hd__o211a_1 _37435_ (.A1(_14553_),
    .A2(_14854_),
    .B1(_14860_),
    .C1(_14859_),
    .X(_14865_));
 sky130_fd_sc_hd__nor2_2 _37436_ (.A(_14864_),
    .B(_14865_),
    .Y(_14866_));
 sky130_fd_sc_hd__nand3_4 _37437_ (.A(_14866_),
    .B(_14790_),
    .C(_14783_),
    .Y(_14867_));
 sky130_fd_sc_hd__nand3_4 _37438_ (.A(_14678_),
    .B(_14863_),
    .C(_14867_),
    .Y(_14868_));
 sky130_fd_sc_hd__nand3_2 _37439_ (.A(_14862_),
    .B(_14790_),
    .C(_14783_),
    .Y(_14869_));
 sky130_fd_sc_hd__nand2_1 _37440_ (.A(_14791_),
    .B(_14866_),
    .Y(_14870_));
 sky130_fd_sc_hd__o2111ai_4 _37441_ (.A1(_14492_),
    .A2(_14579_),
    .B1(_14576_),
    .C1(_14869_),
    .D1(_14870_),
    .Y(_14871_));
 sky130_fd_sc_hd__nand2_1 _37442_ (.A(_14607_),
    .B(_13679_),
    .Y(_14872_));
 sky130_fd_sc_hd__a21oi_4 _37443_ (.A1(_14556_),
    .A2(_14564_),
    .B1(_14568_),
    .Y(_14873_));
 sky130_fd_sc_hd__a21oi_4 _37444_ (.A1(_14539_),
    .A2(_14540_),
    .B1(_14234_),
    .Y(_14874_));
 sky130_fd_sc_hd__nor2_2 _37445_ (.A(_14541_),
    .B(_14874_),
    .Y(_14875_));
 sky130_fd_sc_hd__nand3_4 _37446_ (.A(_14875_),
    .B(_13976_),
    .C(_13977_),
    .Y(_14876_));
 sky130_fd_sc_hd__o211ai_4 _37447_ (.A1(_14541_),
    .A2(_14874_),
    .B1(_13973_),
    .C1(_13970_),
    .Y(_14877_));
 sky130_fd_sc_hd__a21oi_2 _37448_ (.A1(_14876_),
    .A2(_14877_),
    .B1(_14286_),
    .Y(_14878_));
 sky130_fd_sc_hd__and3_1 _37449_ (.A(_14876_),
    .B(_14877_),
    .C(_14278_),
    .X(_14879_));
 sky130_fd_sc_hd__nor2_4 _37450_ (.A(_14535_),
    .B(_14534_),
    .Y(_14880_));
 sky130_fd_sc_hd__nor2_2 _37451_ (.A(_14880_),
    .B(_14548_),
    .Y(_14881_));
 sky130_fd_sc_hd__o21ai_2 _37452_ (.A1(_14878_),
    .A2(_14879_),
    .B1(_14881_),
    .Y(_14882_));
 sky130_fd_sc_hd__nand3_2 _37453_ (.A(_14876_),
    .B(_14877_),
    .C(_14278_),
    .Y(_14883_));
 sky130_fd_sc_hd__a21o_1 _37454_ (.A1(_14876_),
    .A2(_14877_),
    .B1(_14278_),
    .X(_14884_));
 sky130_fd_sc_hd__o211ai_4 _37455_ (.A1(_14880_),
    .A2(_14548_),
    .B1(_14883_),
    .C1(_14884_),
    .Y(_14885_));
 sky130_fd_sc_hd__nand2_1 _37456_ (.A(_14882_),
    .B(_14885_),
    .Y(_14886_));
 sky130_vsdinv _37457_ (.A(_14591_),
    .Y(_14887_));
 sky130_fd_sc_hd__a21oi_4 _37458_ (.A1(_14286_),
    .A2(_14590_),
    .B1(_14887_),
    .Y(_14888_));
 sky130_fd_sc_hd__nand2_4 _37459_ (.A(_14886_),
    .B(_14888_),
    .Y(_14889_));
 sky130_vsdinv _37460_ (.A(_14888_),
    .Y(_14890_));
 sky130_fd_sc_hd__nand3_4 _37461_ (.A(_14882_),
    .B(_14890_),
    .C(_14885_),
    .Y(_14891_));
 sky130_vsdinv _37462_ (.A(_14602_),
    .Y(_14892_));
 sky130_fd_sc_hd__a21oi_2 _37463_ (.A1(_14600_),
    .A2(_14599_),
    .B1(_14598_),
    .Y(_14893_));
 sky130_fd_sc_hd__o21ai_4 _37464_ (.A1(_14892_),
    .A2(_14893_),
    .B1(_14601_),
    .Y(_14894_));
 sky130_fd_sc_hd__a21oi_4 _37465_ (.A1(_14889_),
    .A2(_14891_),
    .B1(_14894_),
    .Y(_14895_));
 sky130_fd_sc_hd__and3_2 _37466_ (.A(_14889_),
    .B(_14894_),
    .C(_14891_),
    .X(_14896_));
 sky130_fd_sc_hd__o21ai_4 _37467_ (.A1(_14895_),
    .A2(_14896_),
    .B1(_14310_),
    .Y(_14897_));
 sky130_fd_sc_hd__a21o_1 _37468_ (.A1(_14889_),
    .A2(_14891_),
    .B1(_14894_),
    .X(_14898_));
 sky130_fd_sc_hd__nand3_4 _37469_ (.A(_14889_),
    .B(_14894_),
    .C(_14891_),
    .Y(_14899_));
 sky130_fd_sc_hd__nand3_4 _37470_ (.A(_14898_),
    .B(_14303_),
    .C(_14899_),
    .Y(_14900_));
 sky130_fd_sc_hd__nand3_4 _37471_ (.A(_14873_),
    .B(_14897_),
    .C(_14900_),
    .Y(_14901_));
 sky130_fd_sc_hd__o21ai_2 _37472_ (.A1(_14895_),
    .A2(_14896_),
    .B1(_13679_),
    .Y(_14902_));
 sky130_fd_sc_hd__o21ai_2 _37473_ (.A1(_14566_),
    .A2(_14567_),
    .B1(_14561_),
    .Y(_14903_));
 sky130_fd_sc_hd__nand3_2 _37474_ (.A(_14898_),
    .B(_14009_),
    .C(_14899_),
    .Y(_14904_));
 sky130_fd_sc_hd__nand3_4 _37475_ (.A(_14902_),
    .B(_14903_),
    .C(_14904_),
    .Y(_14905_));
 sky130_fd_sc_hd__a22oi_4 _37476_ (.A1(_14611_),
    .A2(_14872_),
    .B1(_14901_),
    .B2(_14905_),
    .Y(_14906_));
 sky130_vsdinv _37477_ (.A(_14905_),
    .Y(_14907_));
 sky130_fd_sc_hd__o21ai_2 _37478_ (.A1(_14619_),
    .A2(_14625_),
    .B1(_14901_),
    .Y(_14908_));
 sky130_fd_sc_hd__nor2_2 _37479_ (.A(_14907_),
    .B(_14908_),
    .Y(_14909_));
 sky130_fd_sc_hd__o2bb2ai_4 _37480_ (.A1_N(_14868_),
    .A2_N(_14871_),
    .B1(_14906_),
    .B2(_14909_),
    .Y(_14910_));
 sky130_fd_sc_hd__a32oi_4 _37481_ (.A1(_14873_),
    .A2(_14897_),
    .A3(_14900_),
    .B1(_14607_),
    .B2(_14613_),
    .Y(_14911_));
 sky130_fd_sc_hd__a21oi_4 _37482_ (.A1(_14911_),
    .A2(_14905_),
    .B1(_14906_),
    .Y(_14912_));
 sky130_fd_sc_hd__nand3_4 _37483_ (.A(_14912_),
    .B(_14871_),
    .C(_14868_),
    .Y(_14913_));
 sky130_vsdinv _37484_ (.A(_14585_),
    .Y(_14914_));
 sky130_fd_sc_hd__nand2_1 _37485_ (.A(_14582_),
    .B(_14584_),
    .Y(_14915_));
 sky130_fd_sc_hd__a21oi_2 _37486_ (.A1(_14582_),
    .A2(_14585_),
    .B1(_14584_),
    .Y(_14916_));
 sky130_fd_sc_hd__o22ai_4 _37487_ (.A1(_14914_),
    .A2(_14915_),
    .B1(_14629_),
    .B2(_14916_),
    .Y(_14917_));
 sky130_fd_sc_hd__a21oi_4 _37488_ (.A1(_14910_),
    .A2(_14913_),
    .B1(_14917_),
    .Y(_14918_));
 sky130_fd_sc_hd__and3_1 _37489_ (.A(_14678_),
    .B(_14863_),
    .C(_14867_),
    .X(_14919_));
 sky130_fd_sc_hd__nand2_1 _37490_ (.A(_14912_),
    .B(_14871_),
    .Y(_14920_));
 sky130_fd_sc_hd__o211a_2 _37491_ (.A1(_14919_),
    .A2(_14920_),
    .B1(_14910_),
    .C1(_14917_),
    .X(_14921_));
 sky130_fd_sc_hd__o22ai_4 _37492_ (.A1(_14676_),
    .A2(_14677_),
    .B1(_14918_),
    .B2(_14921_),
    .Y(_14922_));
 sky130_fd_sc_hd__a21o_1 _37493_ (.A1(_14910_),
    .A2(_14913_),
    .B1(_14917_),
    .X(_14923_));
 sky130_fd_sc_hd__nand3_4 _37494_ (.A(_14917_),
    .B(_14910_),
    .C(_14913_),
    .Y(_14924_));
 sky130_fd_sc_hd__nor2_4 _37495_ (.A(_14677_),
    .B(_14676_),
    .Y(_14925_));
 sky130_fd_sc_hd__nand3_2 _37496_ (.A(_14923_),
    .B(_14924_),
    .C(_14925_),
    .Y(_14926_));
 sky130_fd_sc_hd__nand3_4 _37497_ (.A(_14673_),
    .B(_14922_),
    .C(_14926_),
    .Y(_14927_));
 sky130_vsdinv _37498_ (.A(_14674_),
    .Y(_14928_));
 sky130_fd_sc_hd__nor2_4 _37499_ (.A(_14353_),
    .B(_14928_),
    .Y(_14929_));
 sky130_fd_sc_hd__buf_4 _37500_ (.A(_14641_),
    .X(_14930_));
 sky130_fd_sc_hd__buf_6 _37501_ (.A(_14930_),
    .X(_14931_));
 sky130_fd_sc_hd__nor2_2 _37502_ (.A(_14931_),
    .B(_14674_),
    .Y(_14932_));
 sky130_fd_sc_hd__o22ai_4 _37503_ (.A1(_14929_),
    .A2(_14932_),
    .B1(_14918_),
    .B2(_14921_),
    .Y(_14933_));
 sky130_vsdinv _37504_ (.A(_14635_),
    .Y(_14934_));
 sky130_fd_sc_hd__nand2_1 _37505_ (.A(_14648_),
    .B(_14637_),
    .Y(_14935_));
 sky130_fd_sc_hd__o22ai_4 _37506_ (.A1(_14934_),
    .A2(_14935_),
    .B1(_14645_),
    .B2(_14649_),
    .Y(_14936_));
 sky130_fd_sc_hd__o211ai_4 _37507_ (.A1(_14676_),
    .A2(_14677_),
    .B1(_14924_),
    .C1(_14923_),
    .Y(_14937_));
 sky130_fd_sc_hd__nand3_4 _37508_ (.A(_14933_),
    .B(_14936_),
    .C(_14937_),
    .Y(_14938_));
 sky130_fd_sc_hd__clkbuf_4 _37509_ (.A(_14353_),
    .X(_14939_));
 sky130_fd_sc_hd__nor2_4 _37510_ (.A(_14939_),
    .B(_14643_),
    .Y(_14940_));
 sky130_fd_sc_hd__and3_2 _37511_ (.A(_14927_),
    .B(_14938_),
    .C(_14940_),
    .X(_14941_));
 sky130_vsdinv _37512_ (.A(_14647_),
    .Y(_14942_));
 sky130_fd_sc_hd__o21ai_1 _37513_ (.A1(_14343_),
    .A2(_14339_),
    .B1(_14651_),
    .Y(_14943_));
 sky130_fd_sc_hd__o2bb2ai_2 _37514_ (.A1_N(_14333_),
    .A2_N(_14656_),
    .B1(_14942_),
    .B2(_14943_),
    .Y(_14944_));
 sky130_fd_sc_hd__o2bb2ai_1 _37515_ (.A1_N(_14938_),
    .A2_N(_14927_),
    .B1(net412),
    .B2(_14643_),
    .Y(_14945_));
 sky130_fd_sc_hd__nand2_2 _37516_ (.A(_14944_),
    .B(_14945_),
    .Y(_14946_));
 sky130_fd_sc_hd__a21oi_1 _37517_ (.A1(_14927_),
    .A2(_14938_),
    .B1(_14940_),
    .Y(_14947_));
 sky130_fd_sc_hd__o21bai_2 _37518_ (.A1(_14947_),
    .A2(_14941_),
    .B1_N(_14944_),
    .Y(_14948_));
 sky130_fd_sc_hd__o21a_2 _37519_ (.A1(_14941_),
    .A2(_14946_),
    .B1(_14948_),
    .X(_14949_));
 sky130_fd_sc_hd__nand2_2 _37520_ (.A(_14672_),
    .B(_14665_),
    .Y(_14950_));
 sky130_fd_sc_hd__xor2_4 _37521_ (.A(_14949_),
    .B(_14950_),
    .X(_02662_));
 sky130_vsdinv _37522_ (.A(_14938_),
    .Y(_14951_));
 sky130_fd_sc_hd__and2_1 _37523_ (.A(_14927_),
    .B(_14940_),
    .X(_14952_));
 sky130_fd_sc_hd__o21ai_4 _37524_ (.A1(_14925_),
    .A2(_14918_),
    .B1(_14924_),
    .Y(_14953_));
 sky130_fd_sc_hd__o21a_2 _37525_ (.A1(_14709_),
    .A2(_14700_),
    .B1(_14705_),
    .X(_14954_));
 sky130_fd_sc_hd__nand2_2 _37526_ (.A(_11794_),
    .B(_08151_),
    .Y(_14955_));
 sky130_fd_sc_hd__nand2_2 _37527_ (.A(_10989_),
    .B(_08142_),
    .Y(_14956_));
 sky130_fd_sc_hd__nor2_2 _37528_ (.A(_14955_),
    .B(_14956_),
    .Y(_14957_));
 sky130_fd_sc_hd__nand2_2 _37529_ (.A(_09320_),
    .B(_20123_),
    .Y(_14958_));
 sky130_fd_sc_hd__nand2_2 _37530_ (.A(_14955_),
    .B(_14956_),
    .Y(_14959_));
 sky130_fd_sc_hd__nand3b_2 _37531_ (.A_N(_14957_),
    .B(_14958_),
    .C(_14959_),
    .Y(_14960_));
 sky130_vsdinv _37532_ (.A(_14960_),
    .Y(_14961_));
 sky130_fd_sc_hd__and2_1 _37533_ (.A(_14955_),
    .B(_14956_),
    .X(_14962_));
 sky130_vsdinv _37534_ (.A(_14958_),
    .Y(_14963_));
 sky130_fd_sc_hd__o21ai_1 _37535_ (.A1(_14957_),
    .A2(_14962_),
    .B1(_14963_),
    .Y(_14964_));
 sky130_vsdinv _37536_ (.A(_14964_),
    .Y(_14965_));
 sky130_fd_sc_hd__nand3_4 _37537_ (.A(_11778_),
    .B(_11777_),
    .C(_06442_),
    .Y(_14966_));
 sky130_fd_sc_hd__nor2_4 _37538_ (.A(net466),
    .B(_14966_),
    .Y(_14967_));
 sky130_fd_sc_hd__a22oi_4 _37539_ (.A1(_19829_),
    .A2(_07004_),
    .B1(net465),
    .B2(_12487_),
    .Y(_14968_));
 sky130_fd_sc_hd__nand2_4 _37540_ (.A(_10577_),
    .B(_06437_),
    .Y(_14969_));
 sky130_fd_sc_hd__o21ai_4 _37541_ (.A1(_14967_),
    .A2(_14968_),
    .B1(_14969_),
    .Y(_14970_));
 sky130_fd_sc_hd__nand2_1 _37542_ (.A(_10575_),
    .B(_06438_),
    .Y(_14971_));
 sky130_fd_sc_hd__nand3b_4 _37543_ (.A_N(_14971_),
    .B(_18694_),
    .C(_06446_),
    .Y(_14972_));
 sky130_fd_sc_hd__o21ai_2 _37544_ (.A1(net466),
    .A2(_13142_),
    .B1(_14971_),
    .Y(_14973_));
 sky130_vsdinv _37545_ (.A(_14969_),
    .Y(_14974_));
 sky130_fd_sc_hd__nand3_4 _37546_ (.A(_14972_),
    .B(_14973_),
    .C(_14974_),
    .Y(_14975_));
 sky130_fd_sc_hd__o21ai_4 _37547_ (.A1(_14696_),
    .A2(_14691_),
    .B1(_14694_),
    .Y(_14976_));
 sky130_fd_sc_hd__a21oi_4 _37548_ (.A1(_14970_),
    .A2(_14975_),
    .B1(_14976_),
    .Y(_14977_));
 sky130_fd_sc_hd__o21ai_1 _37549_ (.A1(_20139_),
    .A2(_14966_),
    .B1(_14974_),
    .Y(_14978_));
 sky130_fd_sc_hd__o211a_2 _37550_ (.A1(_14968_),
    .A2(_14978_),
    .B1(_14976_),
    .C1(_14970_),
    .X(_14979_));
 sky130_fd_sc_hd__o22ai_4 _37551_ (.A1(_14961_),
    .A2(_14965_),
    .B1(_14977_),
    .B2(_14979_),
    .Y(_14980_));
 sky130_fd_sc_hd__nand2_1 _37552_ (.A(_14970_),
    .B(_14975_),
    .Y(_14981_));
 sky130_fd_sc_hd__a21oi_4 _37553_ (.A1(_14695_),
    .A2(_14697_),
    .B1(_14690_),
    .Y(_14982_));
 sky130_fd_sc_hd__nand2_4 _37554_ (.A(_14981_),
    .B(_14982_),
    .Y(_14983_));
 sky130_fd_sc_hd__nand3_4 _37555_ (.A(_14970_),
    .B(_14976_),
    .C(_14975_),
    .Y(_14984_));
 sky130_fd_sc_hd__o21ai_1 _37556_ (.A1(_14957_),
    .A2(_14962_),
    .B1(_14958_),
    .Y(_14985_));
 sky130_fd_sc_hd__nand3b_1 _37557_ (.A_N(_14957_),
    .B(_14963_),
    .C(_14959_),
    .Y(_14986_));
 sky130_fd_sc_hd__nand2_2 _37558_ (.A(_14985_),
    .B(_14986_),
    .Y(_14987_));
 sky130_fd_sc_hd__nand3_4 _37559_ (.A(_14983_),
    .B(_14984_),
    .C(_14987_),
    .Y(_14988_));
 sky130_fd_sc_hd__nand3_4 _37560_ (.A(_14954_),
    .B(_14980_),
    .C(_14988_),
    .Y(_14989_));
 sky130_fd_sc_hd__o21ai_2 _37561_ (.A1(_14977_),
    .A2(_14979_),
    .B1(_14987_),
    .Y(_14990_));
 sky130_fd_sc_hd__o21ai_4 _37562_ (.A1(_14709_),
    .A2(_14700_),
    .B1(_14705_),
    .Y(_14991_));
 sky130_fd_sc_hd__nand2_2 _37563_ (.A(_14964_),
    .B(_14960_),
    .Y(_14992_));
 sky130_fd_sc_hd__nand3_2 _37564_ (.A(_14983_),
    .B(_14984_),
    .C(_14992_),
    .Y(_14993_));
 sky130_fd_sc_hd__nand3_4 _37565_ (.A(_14990_),
    .B(_14991_),
    .C(_14993_),
    .Y(_14994_));
 sky130_fd_sc_hd__nand2_1 _37566_ (.A(_14989_),
    .B(_14994_),
    .Y(_14995_));
 sky130_fd_sc_hd__o21ai_2 _37567_ (.A1(_14683_),
    .A2(_14684_),
    .B1(_14681_),
    .Y(_14996_));
 sky130_fd_sc_hd__nand2_1 _37568_ (.A(_14683_),
    .B(_14684_),
    .Y(_14997_));
 sky130_fd_sc_hd__nand2_4 _37569_ (.A(_14996_),
    .B(_14997_),
    .Y(_14998_));
 sky130_fd_sc_hd__nand2_2 _37570_ (.A(_11008_),
    .B(_07254_),
    .Y(_14999_));
 sky130_fd_sc_hd__a21o_1 _37571_ (.A1(_11371_),
    .A2(_08060_),
    .B1(_14999_),
    .X(_15000_));
 sky130_fd_sc_hd__nand2_2 _37572_ (.A(_19854_),
    .B(_11487_),
    .Y(_15001_));
 sky130_fd_sc_hd__nand3_2 _37573_ (.A(_14999_),
    .B(_11363_),
    .C(_09921_),
    .Y(_15002_));
 sky130_fd_sc_hd__nand3_4 _37574_ (.A(_15000_),
    .B(_15001_),
    .C(_15002_),
    .Y(_15003_));
 sky130_fd_sc_hd__nand3b_4 _37575_ (.A_N(_14999_),
    .B(_12818_),
    .C(_11062_),
    .Y(_15004_));
 sky130_vsdinv _37576_ (.A(_15001_),
    .Y(_15005_));
 sky130_fd_sc_hd__a22o_1 _37577_ (.A1(_19848_),
    .A2(_12059_),
    .B1(_11371_),
    .B2(_10113_),
    .X(_15006_));
 sky130_fd_sc_hd__nand3_4 _37578_ (.A(_15004_),
    .B(_15005_),
    .C(_15006_),
    .Y(_15007_));
 sky130_fd_sc_hd__nand3b_4 _37579_ (.A_N(_14998_),
    .B(_15003_),
    .C(_15007_),
    .Y(_15008_));
 sky130_vsdinv _37580_ (.A(_10553_),
    .Y(_15009_));
 sky130_fd_sc_hd__buf_2 _37581_ (.A(_15009_),
    .X(_15010_));
 sky130_fd_sc_hd__o31a_2 _37582_ (.A1(_15010_),
    .A2(_10704_),
    .A3(_14716_),
    .B1(_14723_),
    .X(_15011_));
 sky130_fd_sc_hd__a21boi_4 _37583_ (.A1(_15007_),
    .A2(_15003_),
    .B1_N(_14998_),
    .Y(_15012_));
 sky130_fd_sc_hd__nor2_2 _37584_ (.A(_15011_),
    .B(_15012_),
    .Y(_15013_));
 sky130_fd_sc_hd__nand2_1 _37585_ (.A(_15007_),
    .B(_15003_),
    .Y(_15014_));
 sky130_fd_sc_hd__nand2_2 _37586_ (.A(_15014_),
    .B(_14998_),
    .Y(_15015_));
 sky130_fd_sc_hd__nand2_1 _37587_ (.A(_14723_),
    .B(_14720_),
    .Y(_15016_));
 sky130_fd_sc_hd__a21oi_2 _37588_ (.A1(_15015_),
    .A2(_15008_),
    .B1(_15016_),
    .Y(_15017_));
 sky130_fd_sc_hd__a21oi_4 _37589_ (.A1(_15008_),
    .A2(_15013_),
    .B1(_15017_),
    .Y(_15018_));
 sky130_fd_sc_hd__nand2_2 _37590_ (.A(_14995_),
    .B(_15018_),
    .Y(_15019_));
 sky130_fd_sc_hd__a21boi_4 _37591_ (.A1(_14736_),
    .A2(_14711_),
    .B1_N(_14715_),
    .Y(_15020_));
 sky130_fd_sc_hd__nand3b_4 _37592_ (.A_N(_15018_),
    .B(_14989_),
    .C(_14994_),
    .Y(_15021_));
 sky130_fd_sc_hd__nand3_4 _37593_ (.A(_15019_),
    .B(_15020_),
    .C(_15021_),
    .Y(_15022_));
 sky130_fd_sc_hd__a21o_1 _37594_ (.A1(_14989_),
    .A2(_14994_),
    .B1(_15018_),
    .X(_15023_));
 sky130_fd_sc_hd__nand2_1 _37595_ (.A(_14736_),
    .B(_14711_),
    .Y(_15024_));
 sky130_fd_sc_hd__nand2_1 _37596_ (.A(_15024_),
    .B(_14715_),
    .Y(_15025_));
 sky130_fd_sc_hd__nand3_2 _37597_ (.A(_14989_),
    .B(_14994_),
    .C(_15018_),
    .Y(_15026_));
 sky130_fd_sc_hd__nand3_4 _37598_ (.A(_15023_),
    .B(_15025_),
    .C(_15026_),
    .Y(_15027_));
 sky130_vsdinv _37599_ (.A(_14754_),
    .Y(_15028_));
 sky130_fd_sc_hd__and3_1 _37600_ (.A(_14758_),
    .B(_14764_),
    .C(_14766_),
    .X(_15029_));
 sky130_fd_sc_hd__a22oi_4 _37601_ (.A1(_13902_),
    .A2(_10343_),
    .B1(_12447_),
    .B2(_10716_),
    .Y(_15030_));
 sky130_fd_sc_hd__nand3_4 _37602_ (.A(_10916_),
    .B(_07965_),
    .C(_20107_),
    .Y(_15031_));
 sky130_fd_sc_hd__nor2_4 _37603_ (.A(_08037_),
    .B(_15031_),
    .Y(_15032_));
 sky130_fd_sc_hd__nand2_4 _37604_ (.A(_10435_),
    .B(_20101_),
    .Y(_15033_));
 sky130_vsdinv _37605_ (.A(_15033_),
    .Y(_15034_));
 sky130_fd_sc_hd__o21ai_2 _37606_ (.A1(_15030_),
    .A2(_15032_),
    .B1(_15034_),
    .Y(_15035_));
 sky130_fd_sc_hd__a21oi_2 _37607_ (.A1(_14752_),
    .A2(_14749_),
    .B1(_14747_),
    .Y(_15036_));
 sky130_fd_sc_hd__a22o_2 _37608_ (.A1(_13902_),
    .A2(_11723_),
    .B1(_13497_),
    .B2(_10716_),
    .X(_15037_));
 sky130_fd_sc_hd__o211ai_4 _37609_ (.A1(_12100_),
    .A2(_15031_),
    .B1(_15033_),
    .C1(_15037_),
    .Y(_15038_));
 sky130_fd_sc_hd__nand3_4 _37610_ (.A(_15035_),
    .B(_15036_),
    .C(_15038_),
    .Y(_15039_));
 sky130_fd_sc_hd__o21ai_2 _37611_ (.A1(_15030_),
    .A2(_15032_),
    .B1(_15033_),
    .Y(_15040_));
 sky130_fd_sc_hd__o211ai_2 _37612_ (.A1(_08038_),
    .A2(_15031_),
    .B1(_15034_),
    .C1(_15037_),
    .Y(_15041_));
 sky130_fd_sc_hd__o22ai_4 _37613_ (.A1(_09733_),
    .A2(_14746_),
    .B1(_14748_),
    .B2(_14745_),
    .Y(_15042_));
 sky130_fd_sc_hd__nand3_4 _37614_ (.A(_15040_),
    .B(_15041_),
    .C(_15042_),
    .Y(_15043_));
 sky130_fd_sc_hd__nand2_1 _37615_ (.A(_15039_),
    .B(_15043_),
    .Y(_15044_));
 sky130_fd_sc_hd__and4_1 _37616_ (.A(_19870_),
    .B(_07902_),
    .C(_12102_),
    .D(_12103_),
    .X(_15045_));
 sky130_fd_sc_hd__nand2_1 _37617_ (.A(_07479_),
    .B(_09902_),
    .Y(_15046_));
 sky130_fd_sc_hd__a22o_1 _37618_ (.A1(_07483_),
    .A2(_11205_),
    .B1(_10936_),
    .B2(_12109_),
    .X(_15047_));
 sky130_fd_sc_hd__nand3b_2 _37619_ (.A_N(_15045_),
    .B(_15046_),
    .C(_15047_),
    .Y(_15048_));
 sky130_fd_sc_hd__a22oi_2 _37620_ (.A1(_10935_),
    .A2(_11205_),
    .B1(_10945_),
    .B2(_20094_),
    .Y(_15049_));
 sky130_vsdinv _37621_ (.A(_15046_),
    .Y(_15050_));
 sky130_fd_sc_hd__o21ai_1 _37622_ (.A1(_15049_),
    .A2(_15045_),
    .B1(_15050_),
    .Y(_15051_));
 sky130_fd_sc_hd__and2_1 _37623_ (.A(_15048_),
    .B(_15051_),
    .X(_15052_));
 sky130_fd_sc_hd__nand2_2 _37624_ (.A(_15044_),
    .B(_15052_),
    .Y(_15053_));
 sky130_fd_sc_hd__nand2_2 _37625_ (.A(_15048_),
    .B(_15051_),
    .Y(_15054_));
 sky130_fd_sc_hd__nand3_4 _37626_ (.A(_15054_),
    .B(_15039_),
    .C(_15043_),
    .Y(_15055_));
 sky130_fd_sc_hd__a21oi_2 _37627_ (.A1(_14719_),
    .A2(_14723_),
    .B1(_14727_),
    .Y(_15056_));
 sky130_fd_sc_hd__o21ai_4 _37628_ (.A1(_14729_),
    .A2(_15056_),
    .B1(_14728_),
    .Y(_15057_));
 sky130_fd_sc_hd__a21oi_2 _37629_ (.A1(_15053_),
    .A2(_15055_),
    .B1(_15057_),
    .Y(_15058_));
 sky130_vsdinv _37630_ (.A(_14728_),
    .Y(_15059_));
 sky130_fd_sc_hd__o211a_2 _37631_ (.A1(_15059_),
    .A2(_14731_),
    .B1(_15055_),
    .C1(_15053_),
    .X(_15060_));
 sky130_fd_sc_hd__o22ai_2 _37632_ (.A1(_15028_),
    .A2(_15029_),
    .B1(_15058_),
    .B2(_15060_),
    .Y(_15061_));
 sky130_vsdinv _37633_ (.A(_15061_),
    .Y(_15062_));
 sky130_fd_sc_hd__a21o_1 _37634_ (.A1(_15053_),
    .A2(_15055_),
    .B1(_15057_),
    .X(_15063_));
 sky130_fd_sc_hd__nand3_4 _37635_ (.A(_15057_),
    .B(_15055_),
    .C(_15053_),
    .Y(_15064_));
 sky130_fd_sc_hd__nor2_4 _37636_ (.A(_15028_),
    .B(_15029_),
    .Y(_15065_));
 sky130_fd_sc_hd__nand3_2 _37637_ (.A(_15063_),
    .B(_15064_),
    .C(_15065_),
    .Y(_15066_));
 sky130_vsdinv _37638_ (.A(_15066_),
    .Y(_15067_));
 sky130_fd_sc_hd__o2bb2ai_4 _37639_ (.A1_N(_15022_),
    .A2_N(_15027_),
    .B1(_15062_),
    .B2(_15067_),
    .Y(_15068_));
 sky130_fd_sc_hd__o21ai_1 _37640_ (.A1(_15058_),
    .A2(_15060_),
    .B1(_15065_),
    .Y(_15069_));
 sky130_fd_sc_hd__nand3b_1 _37641_ (.A_N(_15065_),
    .B(_15063_),
    .C(_15064_),
    .Y(_15070_));
 sky130_fd_sc_hd__nand2_2 _37642_ (.A(_15069_),
    .B(_15070_),
    .Y(_15071_));
 sky130_fd_sc_hd__nand3_4 _37643_ (.A(_15027_),
    .B(_15022_),
    .C(_15071_),
    .Y(_15072_));
 sky130_fd_sc_hd__a21oi_4 _37644_ (.A1(_14740_),
    .A2(_14743_),
    .B1(_14742_),
    .Y(_15073_));
 sky130_fd_sc_hd__a21o_2 _37645_ (.A1(_14781_),
    .A2(_14744_),
    .B1(_15073_),
    .X(_15074_));
 sky130_fd_sc_hd__a21oi_4 _37646_ (.A1(_15068_),
    .A2(_15072_),
    .B1(_15074_),
    .Y(_15075_));
 sky130_fd_sc_hd__a21oi_2 _37647_ (.A1(_15019_),
    .A2(_15021_),
    .B1(_15020_),
    .Y(_15076_));
 sky130_fd_sc_hd__nand2_1 _37648_ (.A(_15022_),
    .B(_15071_),
    .Y(_15077_));
 sky130_fd_sc_hd__o211a_2 _37649_ (.A1(_15076_),
    .A2(_15077_),
    .B1(_15068_),
    .C1(_15074_),
    .X(_15078_));
 sky130_fd_sc_hd__nand2_2 _37650_ (.A(_06544_),
    .B(_20072_),
    .Y(_15079_));
 sky130_fd_sc_hd__nand2_2 _37651_ (.A(_07422_),
    .B(_10777_),
    .Y(_15080_));
 sky130_fd_sc_hd__nor2_2 _37652_ (.A(_15079_),
    .B(_15080_),
    .Y(_15081_));
 sky130_fd_sc_hd__nand2_4 _37653_ (.A(net503),
    .B(_10700_),
    .Y(_15082_));
 sky130_vsdinv _37654_ (.A(_15082_),
    .Y(_15083_));
 sky130_fd_sc_hd__nand2_2 _37655_ (.A(_15079_),
    .B(_15080_),
    .Y(_15084_));
 sky130_fd_sc_hd__nand3b_4 _37656_ (.A_N(_15081_),
    .B(_15083_),
    .C(_15084_),
    .Y(_15085_));
 sky130_fd_sc_hd__a21o_1 _37657_ (.A1(_06360_),
    .A2(_20069_),
    .B1(_15079_),
    .X(_15086_));
 sky130_fd_sc_hd__a21o_1 _37658_ (.A1(_06358_),
    .A2(_10760_),
    .B1(_15080_),
    .X(_15087_));
 sky130_fd_sc_hd__nand3_4 _37659_ (.A(_15086_),
    .B(_15087_),
    .C(_15082_),
    .Y(_15088_));
 sky130_fd_sc_hd__nor2_1 _37660_ (.A(_14792_),
    .B(_14794_),
    .Y(_15089_));
 sky130_fd_sc_hd__a31o_2 _37661_ (.A1(_14798_),
    .A2(net455),
    .A3(_11604_),
    .B1(_15089_),
    .X(_15090_));
 sky130_fd_sc_hd__a21o_1 _37662_ (.A1(_15085_),
    .A2(_15088_),
    .B1(_15090_),
    .X(_15091_));
 sky130_fd_sc_hd__nand3_4 _37663_ (.A(_15090_),
    .B(_15085_),
    .C(_15088_),
    .Y(_15092_));
 sky130_fd_sc_hd__a21oi_4 _37664_ (.A1(_15091_),
    .A2(_15092_),
    .B1(_14812_),
    .Y(_15093_));
 sky130_fd_sc_hd__and3_2 _37665_ (.A(_15091_),
    .B(_14811_),
    .C(_15092_),
    .X(_15094_));
 sky130_fd_sc_hd__nand2_1 _37666_ (.A(_07294_),
    .B(_20085_),
    .Y(_15095_));
 sky130_fd_sc_hd__a21o_1 _37667_ (.A1(_11094_),
    .A2(_20082_),
    .B1(_15095_),
    .X(_15096_));
 sky130_fd_sc_hd__nand2_1 _37668_ (.A(_07090_),
    .B(_10259_),
    .Y(_15097_));
 sky130_fd_sc_hd__a21o_1 _37669_ (.A1(_11103_),
    .A2(_20086_),
    .B1(_15097_),
    .X(_15098_));
 sky130_fd_sc_hd__o211ai_4 _37670_ (.A1(net443),
    .A2(_12688_),
    .B1(_15096_),
    .C1(_15098_),
    .Y(_15099_));
 sky130_fd_sc_hd__nand3b_4 _37671_ (.A_N(_15095_),
    .B(_11094_),
    .C(_20082_),
    .Y(_15100_));
 sky130_fd_sc_hd__nor2_2 _37672_ (.A(_06528_),
    .B(_11180_),
    .Y(_15101_));
 sky130_fd_sc_hd__nand2_1 _37673_ (.A(_15095_),
    .B(_15097_),
    .Y(_15102_));
 sky130_fd_sc_hd__nand3_4 _37674_ (.A(_15100_),
    .B(_15101_),
    .C(_15102_),
    .Y(_15103_));
 sky130_fd_sc_hd__o21ai_1 _37675_ (.A1(_14759_),
    .A2(_14760_),
    .B1(_14763_),
    .Y(_15104_));
 sky130_fd_sc_hd__nand2_1 _37676_ (.A(_15104_),
    .B(_14765_),
    .Y(_15105_));
 sky130_fd_sc_hd__a21boi_2 _37677_ (.A1(_15099_),
    .A2(_15103_),
    .B1_N(_15105_),
    .Y(_15106_));
 sky130_fd_sc_hd__a21oi_1 _37678_ (.A1(_14759_),
    .A2(_14760_),
    .B1(_14763_),
    .Y(_15107_));
 sky130_fd_sc_hd__o211a_1 _37679_ (.A1(_14761_),
    .A2(_15107_),
    .B1(_15103_),
    .C1(_15099_),
    .X(_15108_));
 sky130_fd_sc_hd__nand2_2 _37680_ (.A(_14825_),
    .B(_14822_),
    .Y(_15109_));
 sky130_fd_sc_hd__o21bai_4 _37681_ (.A1(_15106_),
    .A2(_15108_),
    .B1_N(_15109_),
    .Y(_15110_));
 sky130_fd_sc_hd__nand2_1 _37682_ (.A(_15099_),
    .B(_15103_),
    .Y(_15111_));
 sky130_fd_sc_hd__nand2_2 _37683_ (.A(_15111_),
    .B(_15105_),
    .Y(_15112_));
 sky130_fd_sc_hd__nand3b_4 _37684_ (.A_N(_15105_),
    .B(_15099_),
    .C(_15103_),
    .Y(_15113_));
 sky130_fd_sc_hd__nand3_4 _37685_ (.A(_15112_),
    .B(_15109_),
    .C(_15113_),
    .Y(_15114_));
 sky130_fd_sc_hd__o21ai_4 _37686_ (.A1(_14830_),
    .A2(_14827_),
    .B1(_14833_),
    .Y(_15115_));
 sky130_fd_sc_hd__a21oi_4 _37687_ (.A1(_15110_),
    .A2(_15114_),
    .B1(_15115_),
    .Y(_15116_));
 sky130_fd_sc_hd__nand2_2 _37688_ (.A(_15112_),
    .B(_15109_),
    .Y(_15117_));
 sky130_fd_sc_hd__o211a_2 _37689_ (.A1(_15108_),
    .A2(_15117_),
    .B1(_15115_),
    .C1(_15110_),
    .X(_15118_));
 sky130_fd_sc_hd__o22ai_4 _37690_ (.A1(_15093_),
    .A2(_15094_),
    .B1(_15116_),
    .B2(_15118_),
    .Y(_15119_));
 sky130_fd_sc_hd__a21o_1 _37691_ (.A1(_15110_),
    .A2(_15114_),
    .B1(_15115_),
    .X(_15120_));
 sky130_fd_sc_hd__nor2_4 _37692_ (.A(_15093_),
    .B(_15094_),
    .Y(_15121_));
 sky130_fd_sc_hd__nand3_2 _37693_ (.A(_15110_),
    .B(_15115_),
    .C(_15114_),
    .Y(_15122_));
 sky130_fd_sc_hd__nand3_4 _37694_ (.A(_15120_),
    .B(_15121_),
    .C(_15122_),
    .Y(_15123_));
 sky130_fd_sc_hd__o21ai_4 _37695_ (.A1(_14775_),
    .A2(_14779_),
    .B1(_14772_),
    .Y(_15124_));
 sky130_fd_sc_hd__a21oi_4 _37696_ (.A1(_15119_),
    .A2(_15123_),
    .B1(_15124_),
    .Y(_15125_));
 sky130_vsdinv _37697_ (.A(_14772_),
    .Y(_15126_));
 sky130_fd_sc_hd__o211a_1 _37698_ (.A1(_15126_),
    .A2(_14780_),
    .B1(_15123_),
    .C1(_15119_),
    .X(_15127_));
 sky130_fd_sc_hd__nor2_4 _37699_ (.A(_14846_),
    .B(_14837_),
    .Y(_15128_));
 sky130_fd_sc_hd__nor2_8 _37700_ (.A(_14839_),
    .B(_15128_),
    .Y(_15129_));
 sky130_fd_sc_hd__o21ai_2 _37701_ (.A1(_15125_),
    .A2(_15127_),
    .B1(_15129_),
    .Y(_15130_));
 sky130_fd_sc_hd__a21o_1 _37702_ (.A1(_15119_),
    .A2(_15123_),
    .B1(_15124_),
    .X(_15131_));
 sky130_vsdinv _37703_ (.A(_15129_),
    .Y(_15132_));
 sky130_fd_sc_hd__nand3_4 _37704_ (.A(_15119_),
    .B(_15124_),
    .C(_15123_),
    .Y(_15133_));
 sky130_fd_sc_hd__nand3_2 _37705_ (.A(_15131_),
    .B(_15132_),
    .C(_15133_),
    .Y(_15134_));
 sky130_fd_sc_hd__nand2_4 _37706_ (.A(_15130_),
    .B(_15134_),
    .Y(_15135_));
 sky130_fd_sc_hd__o21ai_2 _37707_ (.A1(_15075_),
    .A2(_15078_),
    .B1(_15135_),
    .Y(_15136_));
 sky130_fd_sc_hd__o21ai_1 _37708_ (.A1(_15125_),
    .A2(_15127_),
    .B1(_15132_),
    .Y(_15137_));
 sky130_fd_sc_hd__nand3_2 _37709_ (.A(_15131_),
    .B(_15133_),
    .C(_15129_),
    .Y(_15138_));
 sky130_fd_sc_hd__nand2_1 _37710_ (.A(_15068_),
    .B(_15072_),
    .Y(_15139_));
 sky130_fd_sc_hd__a21oi_4 _37711_ (.A1(_14781_),
    .A2(_14744_),
    .B1(_15073_),
    .Y(_15140_));
 sky130_fd_sc_hd__a22oi_2 _37712_ (.A1(_15137_),
    .A2(_15138_),
    .B1(_15139_),
    .B2(_15140_),
    .Y(_15141_));
 sky130_fd_sc_hd__nand3_2 _37713_ (.A(_15074_),
    .B(_15072_),
    .C(_15068_),
    .Y(_15142_));
 sky130_fd_sc_hd__nand2_1 _37714_ (.A(_15141_),
    .B(_15142_),
    .Y(_15143_));
 sky130_fd_sc_hd__a21oi_4 _37715_ (.A1(_14786_),
    .A2(_14789_),
    .B1(_14788_),
    .Y(_15144_));
 sky130_fd_sc_hd__a31o_1 _37716_ (.A1(_14790_),
    .A2(_14861_),
    .A3(_14856_),
    .B1(_15144_),
    .X(_15145_));
 sky130_fd_sc_hd__nand3_4 _37717_ (.A(_15136_),
    .B(_15143_),
    .C(_15145_),
    .Y(_15146_));
 sky130_vsdinv _37718_ (.A(_15138_),
    .Y(_15147_));
 sky130_vsdinv _37719_ (.A(_15137_),
    .Y(_15148_));
 sky130_fd_sc_hd__o22ai_4 _37720_ (.A1(_15147_),
    .A2(_15148_),
    .B1(_15075_),
    .B2(_15078_),
    .Y(_15149_));
 sky130_fd_sc_hd__a31oi_4 _37721_ (.A1(_14790_),
    .A2(_14861_),
    .A3(_14856_),
    .B1(_15144_),
    .Y(_15150_));
 sky130_fd_sc_hd__nand2_2 _37722_ (.A(_15139_),
    .B(_15140_),
    .Y(_15151_));
 sky130_fd_sc_hd__nand3_2 _37723_ (.A(_15151_),
    .B(_15142_),
    .C(_15135_),
    .Y(_15152_));
 sky130_fd_sc_hd__nand3_4 _37724_ (.A(_15149_),
    .B(_15150_),
    .C(_15152_),
    .Y(_15153_));
 sky130_fd_sc_hd__nand2_1 _37725_ (.A(_15146_),
    .B(_15153_),
    .Y(_15154_));
 sky130_fd_sc_hd__a21oi_4 _37726_ (.A1(_14857_),
    .A2(_14859_),
    .B1(_14853_),
    .Y(_15155_));
 sky130_fd_sc_hd__o21ai_2 _37727_ (.A1(_06344_),
    .A2(_06909_),
    .B1(_12348_),
    .Y(_15156_));
 sky130_fd_sc_hd__o21a_2 _37728_ (.A1(_05632_),
    .A2(_15156_),
    .B1(_14808_),
    .X(_15157_));
 sky130_fd_sc_hd__nand3_4 _37729_ (.A(_13976_),
    .B(_15157_),
    .C(_13977_),
    .Y(_15158_));
 sky130_fd_sc_hd__o21ai_4 _37730_ (.A1(_05633_),
    .A2(_15156_),
    .B1(_14808_),
    .Y(_15159_));
 sky130_fd_sc_hd__nand3_4 _37731_ (.A(_13970_),
    .B(_13973_),
    .C(_15159_),
    .Y(_15160_));
 sky130_fd_sc_hd__nand2_1 _37732_ (.A(_15158_),
    .B(_15160_),
    .Y(_15161_));
 sky130_fd_sc_hd__nor2_4 _37733_ (.A(_13969_),
    .B(_13971_),
    .Y(_15162_));
 sky130_fd_sc_hd__nand2_4 _37734_ (.A(_15161_),
    .B(_15162_),
    .Y(_15163_));
 sky130_fd_sc_hd__nand3_4 _37735_ (.A(_15158_),
    .B(_15160_),
    .C(_14278_),
    .Y(_15164_));
 sky130_fd_sc_hd__nand2_2 _37736_ (.A(_15163_),
    .B(_15164_),
    .Y(_15165_));
 sky130_fd_sc_hd__a21oi_2 _37737_ (.A1(_14803_),
    .A2(_14811_),
    .B1(_14842_),
    .Y(_15166_));
 sky130_fd_sc_hd__nand2_2 _37738_ (.A(_15165_),
    .B(_15166_),
    .Y(_15167_));
 sky130_fd_sc_hd__o21ai_4 _37739_ (.A1(_14843_),
    .A2(_14841_),
    .B1(_14805_),
    .Y(_15168_));
 sky130_fd_sc_hd__nand3_4 _37740_ (.A(_15168_),
    .B(_15164_),
    .C(_15163_),
    .Y(_15169_));
 sky130_vsdinv _37741_ (.A(_14877_),
    .Y(_15170_));
 sky130_fd_sc_hd__a21oi_4 _37742_ (.A1(_14286_),
    .A2(_14876_),
    .B1(_15170_),
    .Y(_15171_));
 sky130_vsdinv _37743_ (.A(_15171_),
    .Y(_15172_));
 sky130_fd_sc_hd__a21oi_4 _37744_ (.A1(_15167_),
    .A2(_15169_),
    .B1(_15172_),
    .Y(_15173_));
 sky130_fd_sc_hd__and3_1 _37745_ (.A(_15167_),
    .B(_15172_),
    .C(_15169_),
    .X(_15174_));
 sky130_fd_sc_hd__o31a_1 _37746_ (.A1(_14878_),
    .A2(_14881_),
    .A3(_14879_),
    .B1(_14891_),
    .X(_15175_));
 sky130_fd_sc_hd__o21ai_4 _37747_ (.A1(_15173_),
    .A2(_15174_),
    .B1(_15175_),
    .Y(_15176_));
 sky130_fd_sc_hd__nand3_2 _37748_ (.A(_15167_),
    .B(_15169_),
    .C(_15172_),
    .Y(_15177_));
 sky130_fd_sc_hd__nand2_2 _37749_ (.A(_14891_),
    .B(_14885_),
    .Y(_15178_));
 sky130_fd_sc_hd__nand3b_4 _37750_ (.A_N(_15173_),
    .B(_15177_),
    .C(_15178_),
    .Y(_15179_));
 sky130_fd_sc_hd__nand2_1 _37751_ (.A(_15176_),
    .B(_15179_),
    .Y(_15180_));
 sky130_fd_sc_hd__nand2_1 _37752_ (.A(_15180_),
    .B(_14310_),
    .Y(_15181_));
 sky130_fd_sc_hd__nand3_2 _37753_ (.A(_15176_),
    .B(_15179_),
    .C(_14303_),
    .Y(_15182_));
 sky130_fd_sc_hd__nand3_4 _37754_ (.A(_15155_),
    .B(_15181_),
    .C(_15182_),
    .Y(_15183_));
 sky130_fd_sc_hd__o21ai_2 _37755_ (.A1(_14855_),
    .A2(_14851_),
    .B1(_14860_),
    .Y(_15184_));
 sky130_fd_sc_hd__o2bb2ai_1 _37756_ (.A1_N(_15179_),
    .A2_N(_15176_),
    .B1(_13689_),
    .B2(_13675_),
    .Y(_15185_));
 sky130_fd_sc_hd__nand3_2 _37757_ (.A(_15176_),
    .B(_15179_),
    .C(_13686_),
    .Y(_15186_));
 sky130_fd_sc_hd__nand3_4 _37758_ (.A(_15184_),
    .B(_15185_),
    .C(_15186_),
    .Y(_15187_));
 sky130_fd_sc_hd__nor2_1 _37759_ (.A(_14303_),
    .B(_14895_),
    .Y(_15188_));
 sky130_fd_sc_hd__or2_1 _37760_ (.A(_14896_),
    .B(_15188_),
    .X(_15189_));
 sky130_fd_sc_hd__a21oi_2 _37761_ (.A1(_15183_),
    .A2(_15187_),
    .B1(_15189_),
    .Y(_15190_));
 sky130_fd_sc_hd__o211a_1 _37762_ (.A1(_14896_),
    .A2(_15188_),
    .B1(_15187_),
    .C1(_15183_),
    .X(_15191_));
 sky130_fd_sc_hd__nor2_2 _37763_ (.A(_15190_),
    .B(_15191_),
    .Y(_15192_));
 sky130_fd_sc_hd__nand2_1 _37764_ (.A(_15154_),
    .B(_15192_),
    .Y(_15193_));
 sky130_fd_sc_hd__a21oi_4 _37765_ (.A1(_14912_),
    .A2(_14871_),
    .B1(_14919_),
    .Y(_15194_));
 sky130_fd_sc_hd__nand3_1 _37766_ (.A(_15189_),
    .B(_15183_),
    .C(_15187_),
    .Y(_15195_));
 sky130_fd_sc_hd__or2b_1 _37767_ (.A(_15190_),
    .B_N(_15195_),
    .X(_15196_));
 sky130_fd_sc_hd__nand3_2 _37768_ (.A(_15196_),
    .B(_15153_),
    .C(_15146_),
    .Y(_15197_));
 sky130_fd_sc_hd__nand3_4 _37769_ (.A(_15193_),
    .B(_15194_),
    .C(_15197_),
    .Y(_15198_));
 sky130_fd_sc_hd__nand2_1 _37770_ (.A(_15154_),
    .B(_15196_),
    .Y(_15199_));
 sky130_fd_sc_hd__nand2_1 _37771_ (.A(_14920_),
    .B(_14868_),
    .Y(_15200_));
 sky130_fd_sc_hd__nand3_2 _37772_ (.A(_15192_),
    .B(_15146_),
    .C(_15153_),
    .Y(_15201_));
 sky130_fd_sc_hd__nand3_4 _37773_ (.A(_15199_),
    .B(_15200_),
    .C(_15201_),
    .Y(_15202_));
 sky130_fd_sc_hd__nand2_4 _37774_ (.A(_14908_),
    .B(_14905_),
    .Y(_15203_));
 sky130_fd_sc_hd__nor2_8 _37775_ (.A(_14641_),
    .B(_15203_),
    .Y(_15204_));
 sky130_vsdinv _37776_ (.A(_15203_),
    .Y(_15205_));
 sky130_fd_sc_hd__nor2_8 _37777_ (.A(_13739_),
    .B(_15205_),
    .Y(_15206_));
 sky130_fd_sc_hd__nor2_8 _37778_ (.A(_15204_),
    .B(_15206_),
    .Y(_15207_));
 sky130_vsdinv _37779_ (.A(_15207_),
    .Y(_15208_));
 sky130_fd_sc_hd__a21o_1 _37780_ (.A1(_15198_),
    .A2(_15202_),
    .B1(_15208_),
    .X(_15209_));
 sky130_fd_sc_hd__nand3_2 _37781_ (.A(_15208_),
    .B(_15198_),
    .C(_15202_),
    .Y(_15210_));
 sky130_fd_sc_hd__nand3b_4 _37782_ (.A_N(_14953_),
    .B(_15209_),
    .C(_15210_),
    .Y(_15211_));
 sky130_fd_sc_hd__o2bb2ai_4 _37783_ (.A1_N(_15202_),
    .A2_N(_15198_),
    .B1(_15206_),
    .B2(_15204_),
    .Y(_15212_));
 sky130_fd_sc_hd__nand3_4 _37784_ (.A(_15198_),
    .B(_15202_),
    .C(_15207_),
    .Y(_15213_));
 sky130_fd_sc_hd__nand3_4 _37785_ (.A(_15212_),
    .B(_15213_),
    .C(_14953_),
    .Y(_15214_));
 sky130_fd_sc_hd__nand3_2 _37786_ (.A(_15211_),
    .B(_14929_),
    .C(_15214_),
    .Y(_15215_));
 sky130_fd_sc_hd__nand2_1 _37787_ (.A(_15211_),
    .B(_15214_),
    .Y(_15216_));
 sky130_vsdinv _37788_ (.A(_14929_),
    .Y(_15217_));
 sky130_fd_sc_hd__nand2_1 _37789_ (.A(_15216_),
    .B(_15217_),
    .Y(_15218_));
 sky130_fd_sc_hd__o211ai_4 _37790_ (.A1(_14951_),
    .A2(_14952_),
    .B1(_15215_),
    .C1(_15218_),
    .Y(_15219_));
 sky130_fd_sc_hd__nand2_1 _37791_ (.A(_15216_),
    .B(_14929_),
    .Y(_15220_));
 sky130_fd_sc_hd__a21oi_2 _37792_ (.A1(_14927_),
    .A2(_14940_),
    .B1(_14951_),
    .Y(_15221_));
 sky130_fd_sc_hd__nand3_2 _37793_ (.A(_15211_),
    .B(_15217_),
    .C(_15214_),
    .Y(_15222_));
 sky130_fd_sc_hd__nand3_4 _37794_ (.A(_15220_),
    .B(_15221_),
    .C(_15222_),
    .Y(_15223_));
 sky130_fd_sc_hd__nand2_1 _37795_ (.A(_15219_),
    .B(_15223_),
    .Y(_15224_));
 sky130_vsdinv _37796_ (.A(_15224_),
    .Y(_15225_));
 sky130_fd_sc_hd__o2111ai_4 _37797_ (.A1(_14941_),
    .A2(_14946_),
    .B1(_14665_),
    .C1(_14948_),
    .D1(_14660_),
    .Y(_15226_));
 sky130_fd_sc_hd__and2_1 _37798_ (.A(_14047_),
    .B(_14048_),
    .X(_15227_));
 sky130_fd_sc_hd__nand3b_4 _37799_ (.A_N(_15226_),
    .B(_15227_),
    .C(_14360_),
    .Y(_15228_));
 sky130_fd_sc_hd__nand3_1 _37800_ (.A(_14927_),
    .B(_14938_),
    .C(_14940_),
    .Y(_15229_));
 sky130_fd_sc_hd__a21oi_1 _37801_ (.A1(_14945_),
    .A2(_15229_),
    .B1(_14944_),
    .Y(_15230_));
 sky130_fd_sc_hd__o22ai_1 _37802_ (.A1(_14941_),
    .A2(_14946_),
    .B1(_15230_),
    .B2(_14665_),
    .Y(_15231_));
 sky130_fd_sc_hd__o21bai_1 _37803_ (.A1(_15226_),
    .A2(_14669_),
    .B1_N(_15231_),
    .Y(_15232_));
 sky130_fd_sc_hd__o21bai_4 _37804_ (.A1(_15228_),
    .A2(_14056_),
    .B1_N(_15232_),
    .Y(_15233_));
 sky130_fd_sc_hd__xor2_4 _37805_ (.A(_15225_),
    .B(_15233_),
    .X(_02663_));
 sky130_fd_sc_hd__and2_1 _37806_ (.A(_15133_),
    .B(_15129_),
    .X(_15234_));
 sky130_fd_sc_hd__a21oi_4 _37807_ (.A1(_15158_),
    .A2(_15160_),
    .B1(_14286_),
    .Y(_15235_));
 sky130_vsdinv _37808_ (.A(_15164_),
    .Y(_15236_));
 sky130_fd_sc_hd__a21oi_2 _37809_ (.A1(_15085_),
    .A2(_15088_),
    .B1(_15090_),
    .Y(_15237_));
 sky130_fd_sc_hd__o21a_1 _37810_ (.A1(_14843_),
    .A2(_15237_),
    .B1(_15092_),
    .X(_15238_));
 sky130_fd_sc_hd__o21ai_4 _37811_ (.A1(_15235_),
    .A2(_15236_),
    .B1(_15238_),
    .Y(_15239_));
 sky130_fd_sc_hd__o21ai_2 _37812_ (.A1(_14844_),
    .A2(_15237_),
    .B1(_15092_),
    .Y(_15240_));
 sky130_fd_sc_hd__nand3_4 _37813_ (.A(_15240_),
    .B(_15164_),
    .C(_15163_),
    .Y(_15241_));
 sky130_vsdinv _37814_ (.A(_15160_),
    .Y(_15242_));
 sky130_fd_sc_hd__and2_1 _37815_ (.A(_15158_),
    .B(_14278_),
    .X(_15243_));
 sky130_fd_sc_hd__or2_4 _37816_ (.A(_15242_),
    .B(_15243_),
    .X(_15244_));
 sky130_fd_sc_hd__a21oi_4 _37817_ (.A1(_15239_),
    .A2(_15241_),
    .B1(_15244_),
    .Y(_15245_));
 sky130_fd_sc_hd__o211a_1 _37818_ (.A1(_15242_),
    .A2(_15243_),
    .B1(_15241_),
    .C1(_15239_),
    .X(_15246_));
 sky130_vsdinv _37819_ (.A(_15169_),
    .Y(_15247_));
 sky130_fd_sc_hd__a21oi_2 _37820_ (.A1(_15163_),
    .A2(_15164_),
    .B1(_15168_),
    .Y(_15248_));
 sky130_fd_sc_hd__nor2_4 _37821_ (.A(_15171_),
    .B(_15248_),
    .Y(_15249_));
 sky130_fd_sc_hd__nor2_2 _37822_ (.A(_15247_),
    .B(_15249_),
    .Y(_15250_));
 sky130_fd_sc_hd__o21ai_4 _37823_ (.A1(_15245_),
    .A2(_15246_),
    .B1(_15250_),
    .Y(_15251_));
 sky130_fd_sc_hd__nand3_4 _37824_ (.A(_15244_),
    .B(_15239_),
    .C(_15241_),
    .Y(_15252_));
 sky130_fd_sc_hd__nand2_1 _37825_ (.A(_15239_),
    .B(_15241_),
    .Y(_15253_));
 sky130_fd_sc_hd__nor2_1 _37826_ (.A(_15242_),
    .B(_15243_),
    .Y(_15254_));
 sky130_fd_sc_hd__nand2_1 _37827_ (.A(_15253_),
    .B(_15254_),
    .Y(_15255_));
 sky130_fd_sc_hd__o211ai_4 _37828_ (.A1(_15247_),
    .A2(_15249_),
    .B1(_15252_),
    .C1(_15255_),
    .Y(_15256_));
 sky130_fd_sc_hd__a22oi_4 _37829_ (.A1(_13964_),
    .A2(_13965_),
    .B1(_15251_),
    .B2(_15256_),
    .Y(_15257_));
 sky130_fd_sc_hd__o2bb2ai_1 _37830_ (.A1_N(_15253_),
    .A2_N(_15254_),
    .B1(_15247_),
    .B2(_15249_),
    .Y(_15258_));
 sky130_fd_sc_hd__o211a_1 _37831_ (.A1(_15246_),
    .A2(_15258_),
    .B1(_13686_),
    .C1(_15251_),
    .X(_15259_));
 sky130_fd_sc_hd__o22ai_4 _37832_ (.A1(_15125_),
    .A2(_15234_),
    .B1(_15257_),
    .B2(_15259_),
    .Y(_15260_));
 sky130_vsdinv _37833_ (.A(_15256_),
    .Y(_15261_));
 sky130_fd_sc_hd__nand2_2 _37834_ (.A(_15251_),
    .B(_13686_),
    .Y(_15262_));
 sky130_fd_sc_hd__o21ai_2 _37835_ (.A1(_15129_),
    .A2(_15125_),
    .B1(_15133_),
    .Y(_15263_));
 sky130_fd_sc_hd__a21o_1 _37836_ (.A1(_15251_),
    .A2(_15256_),
    .B1(_13686_),
    .X(_15264_));
 sky130_fd_sc_hd__o211ai_4 _37837_ (.A1(_15261_),
    .A2(_15262_),
    .B1(_15263_),
    .C1(_15264_),
    .Y(_15265_));
 sky130_fd_sc_hd__a21bo_2 _37838_ (.A1(_14009_),
    .A2(_15176_),
    .B1_N(_15179_),
    .X(_15266_));
 sky130_fd_sc_hd__a21oi_4 _37839_ (.A1(_15260_),
    .A2(_15265_),
    .B1(_15266_),
    .Y(_15267_));
 sky130_fd_sc_hd__and3_2 _37840_ (.A(_15260_),
    .B(_15265_),
    .C(_15266_),
    .X(_15268_));
 sky130_fd_sc_hd__nand2_1 _37841_ (.A(_15135_),
    .B(_15142_),
    .Y(_15269_));
 sky130_fd_sc_hd__nand2_2 _37842_ (.A(_07088_),
    .B(_20081_),
    .Y(_15270_));
 sky130_fd_sc_hd__nand2_2 _37843_ (.A(_07291_),
    .B(_10256_),
    .Y(_15271_));
 sky130_fd_sc_hd__nor2_2 _37844_ (.A(_15270_),
    .B(_15271_),
    .Y(_15272_));
 sky130_fd_sc_hd__and2_1 _37845_ (.A(_15270_),
    .B(_15271_),
    .X(_15273_));
 sky130_fd_sc_hd__nor2_2 _37846_ (.A(net443),
    .B(_10772_),
    .Y(_15274_));
 sky130_fd_sc_hd__o21bai_4 _37847_ (.A1(_15272_),
    .A2(_15273_),
    .B1_N(_15274_),
    .Y(_15275_));
 sky130_fd_sc_hd__or2_2 _37848_ (.A(_15270_),
    .B(_15271_),
    .X(_15276_));
 sky130_fd_sc_hd__nand2_1 _37849_ (.A(_15270_),
    .B(_15271_),
    .Y(_15277_));
 sky130_fd_sc_hd__nand3_4 _37850_ (.A(_15276_),
    .B(_15274_),
    .C(_15277_),
    .Y(_15278_));
 sky130_fd_sc_hd__a21o_2 _37851_ (.A1(_15047_),
    .A2(_15050_),
    .B1(_15045_),
    .X(_15279_));
 sky130_fd_sc_hd__a21oi_4 _37852_ (.A1(_15275_),
    .A2(_15278_),
    .B1(_15279_),
    .Y(_15280_));
 sky130_fd_sc_hd__nor2_1 _37853_ (.A(_15046_),
    .B(_15049_),
    .Y(_15281_));
 sky130_fd_sc_hd__o211a_1 _37854_ (.A1(_15045_),
    .A2(_15281_),
    .B1(_15278_),
    .C1(_15275_),
    .X(_15282_));
 sky130_fd_sc_hd__nand2_2 _37855_ (.A(_15103_),
    .B(_15100_),
    .Y(_15283_));
 sky130_vsdinv _37856_ (.A(_15283_),
    .Y(_15284_));
 sky130_fd_sc_hd__o21ai_4 _37857_ (.A1(_15280_),
    .A2(_15282_),
    .B1(_15284_),
    .Y(_15285_));
 sky130_fd_sc_hd__a21o_1 _37858_ (.A1(_15275_),
    .A2(_15278_),
    .B1(_15279_),
    .X(_15286_));
 sky130_fd_sc_hd__nand3_4 _37859_ (.A(_15275_),
    .B(_15278_),
    .C(_15279_),
    .Y(_15287_));
 sky130_fd_sc_hd__nand3_4 _37860_ (.A(_15286_),
    .B(_15283_),
    .C(_15287_),
    .Y(_15288_));
 sky130_fd_sc_hd__nand2_4 _37861_ (.A(_15117_),
    .B(_15113_),
    .Y(_15289_));
 sky130_fd_sc_hd__a21oi_4 _37862_ (.A1(_15285_),
    .A2(_15288_),
    .B1(_15289_),
    .Y(_15290_));
 sky130_fd_sc_hd__and3_2 _37863_ (.A(_15285_),
    .B(_15289_),
    .C(_15288_),
    .X(_15291_));
 sky130_fd_sc_hd__nand2_2 _37864_ (.A(_06544_),
    .B(_10777_),
    .Y(_15292_));
 sky130_fd_sc_hd__nand2_2 _37865_ (.A(_14806_),
    .B(_06359_),
    .Y(_15293_));
 sky130_fd_sc_hd__o21ai_1 _37866_ (.A1(_15292_),
    .A2(_15293_),
    .B1(_15082_),
    .Y(_15294_));
 sky130_fd_sc_hd__a21o_1 _37867_ (.A1(_15292_),
    .A2(_15293_),
    .B1(_15294_),
    .X(_15295_));
 sky130_fd_sc_hd__nor2_1 _37868_ (.A(_15292_),
    .B(_15293_),
    .Y(_15296_));
 sky130_fd_sc_hd__and2_1 _37869_ (.A(_15292_),
    .B(_15293_),
    .X(_15297_));
 sky130_fd_sc_hd__o21ai_2 _37870_ (.A1(_15296_),
    .A2(_15297_),
    .B1(_15083_),
    .Y(_15298_));
 sky130_fd_sc_hd__a21oi_4 _37871_ (.A1(_15083_),
    .A2(_15084_),
    .B1(_15081_),
    .Y(_15299_));
 sky130_fd_sc_hd__a21o_2 _37872_ (.A1(_15295_),
    .A2(_15298_),
    .B1(_15299_),
    .X(_15300_));
 sky130_vsdinv _37873_ (.A(_15300_),
    .Y(_15301_));
 sky130_fd_sc_hd__nand3_4 _37874_ (.A(_15295_),
    .B(_15298_),
    .C(_15299_),
    .Y(_15302_));
 sky130_fd_sc_hd__nand2_4 _37875_ (.A(_15302_),
    .B(_14811_),
    .Y(_15303_));
 sky130_fd_sc_hd__a21o_1 _37876_ (.A1(_15300_),
    .A2(_15302_),
    .B1(_14811_),
    .X(_15304_));
 sky130_fd_sc_hd__o21ai_4 _37877_ (.A1(_15301_),
    .A2(_15303_),
    .B1(_15304_),
    .Y(_15305_));
 sky130_fd_sc_hd__o21ai_2 _37878_ (.A1(_15290_),
    .A2(_15291_),
    .B1(_15305_),
    .Y(_15306_));
 sky130_fd_sc_hd__nand2_2 _37879_ (.A(_15066_),
    .B(_15064_),
    .Y(_15307_));
 sky130_fd_sc_hd__a21o_2 _37880_ (.A1(_15285_),
    .A2(_15288_),
    .B1(_15289_),
    .X(_15308_));
 sky130_fd_sc_hd__nand3_4 _37881_ (.A(_15285_),
    .B(_15289_),
    .C(_15288_),
    .Y(_15309_));
 sky130_fd_sc_hd__nand3b_4 _37882_ (.A_N(_15305_),
    .B(_15308_),
    .C(_15309_),
    .Y(_15310_));
 sky130_fd_sc_hd__nand3_4 _37883_ (.A(_15306_),
    .B(_15307_),
    .C(_15310_),
    .Y(_15311_));
 sky130_fd_sc_hd__o21bai_4 _37884_ (.A1(_15290_),
    .A2(_15291_),
    .B1_N(_15305_),
    .Y(_15312_));
 sky130_fd_sc_hd__a21oi_4 _37885_ (.A1(_15063_),
    .A2(_15065_),
    .B1(_15060_),
    .Y(_15313_));
 sky130_fd_sc_hd__nand3_4 _37886_ (.A(_15308_),
    .B(_15305_),
    .C(_15309_),
    .Y(_15314_));
 sky130_fd_sc_hd__nand3_4 _37887_ (.A(_15312_),
    .B(_15313_),
    .C(_15314_),
    .Y(_15315_));
 sky130_fd_sc_hd__nor2_2 _37888_ (.A(_15121_),
    .B(_15118_),
    .Y(_15316_));
 sky130_fd_sc_hd__nor2_4 _37889_ (.A(_15116_),
    .B(_15316_),
    .Y(_15317_));
 sky130_fd_sc_hd__a21oi_2 _37890_ (.A1(_15311_),
    .A2(_15315_),
    .B1(_15317_),
    .Y(_15318_));
 sky130_fd_sc_hd__nand3_1 _37891_ (.A(_15311_),
    .B(_15315_),
    .C(_15317_),
    .Y(_15319_));
 sky130_vsdinv _37892_ (.A(_15319_),
    .Y(_15320_));
 sky130_vsdinv _37893_ (.A(_14975_),
    .Y(_15321_));
 sky130_fd_sc_hd__nand2_1 _37894_ (.A(_14970_),
    .B(_14976_),
    .Y(_15322_));
 sky130_fd_sc_hd__a2bb2oi_4 _37895_ (.A1_N(_15321_),
    .A2_N(_15322_),
    .B1(_14992_),
    .B2(_14983_),
    .Y(_15323_));
 sky130_fd_sc_hd__nand2_4 _37896_ (.A(_19835_),
    .B(_07709_),
    .Y(_15324_));
 sky130_fd_sc_hd__nand2_4 _37897_ (.A(_10989_),
    .B(_07567_),
    .Y(_15325_));
 sky130_fd_sc_hd__nor2_4 _37898_ (.A(_15324_),
    .B(_15325_),
    .Y(_15326_));
 sky130_fd_sc_hd__nand2_2 _37899_ (.A(_15324_),
    .B(_15325_),
    .Y(_15327_));
 sky130_vsdinv _37900_ (.A(_15327_),
    .Y(_15328_));
 sky130_fd_sc_hd__nand2_2 _37901_ (.A(_19844_),
    .B(_11061_),
    .Y(_15329_));
 sky130_vsdinv _37902_ (.A(_15329_),
    .Y(_15330_));
 sky130_fd_sc_hd__o21a_1 _37903_ (.A1(_15326_),
    .A2(_15328_),
    .B1(_15330_),
    .X(_15331_));
 sky130_vsdinv _37904_ (.A(_15326_),
    .Y(_15332_));
 sky130_fd_sc_hd__nand3_2 _37905_ (.A(_15332_),
    .B(_15329_),
    .C(_15327_),
    .Y(_15333_));
 sky130_vsdinv _37906_ (.A(_15333_),
    .Y(_15334_));
 sky130_fd_sc_hd__nand3_4 _37907_ (.A(_10973_),
    .B(_11783_),
    .C(_07003_),
    .Y(_15335_));
 sky130_fd_sc_hd__nor2_4 _37908_ (.A(_20136_),
    .B(_15335_),
    .Y(_15336_));
 sky130_fd_sc_hd__a22oi_4 _37909_ (.A1(_12492_),
    .A2(_10941_),
    .B1(_06722_),
    .B2(_13139_),
    .Y(_15337_));
 sky130_fd_sc_hd__nand2_4 _37910_ (.A(_10573_),
    .B(_06714_),
    .Y(_15338_));
 sky130_fd_sc_hd__o21ai_4 _37911_ (.A1(_15336_),
    .A2(_15337_),
    .B1(_15338_),
    .Y(_15339_));
 sky130_fd_sc_hd__nand2_2 _37912_ (.A(_11783_),
    .B(_20133_),
    .Y(_15340_));
 sky130_fd_sc_hd__nand3b_4 _37913_ (.A_N(_15340_),
    .B(_18694_),
    .C(_07510_),
    .Y(_15341_));
 sky130_fd_sc_hd__o21ai_4 _37914_ (.A1(_06312_),
    .A2(_13142_),
    .B1(_15340_),
    .Y(_15342_));
 sky130_vsdinv _37915_ (.A(_15338_),
    .Y(_15343_));
 sky130_fd_sc_hd__nand3_4 _37916_ (.A(_15341_),
    .B(_15342_),
    .C(_15343_),
    .Y(_15344_));
 sky130_fd_sc_hd__o21ai_4 _37917_ (.A1(_14969_),
    .A2(_14968_),
    .B1(_14972_),
    .Y(_15345_));
 sky130_fd_sc_hd__a21oi_4 _37918_ (.A1(_15339_),
    .A2(_15344_),
    .B1(_15345_),
    .Y(_15346_));
 sky130_fd_sc_hd__o21ai_1 _37919_ (.A1(_20136_),
    .A2(_15335_),
    .B1(_15343_),
    .Y(_15347_));
 sky130_fd_sc_hd__o211a_2 _37920_ (.A1(_15337_),
    .A2(_15347_),
    .B1(_15345_),
    .C1(_15339_),
    .X(_15348_));
 sky130_fd_sc_hd__o22ai_4 _37921_ (.A1(_15331_),
    .A2(_15334_),
    .B1(_15346_),
    .B2(_15348_),
    .Y(_15349_));
 sky130_fd_sc_hd__nand2_1 _37922_ (.A(_15339_),
    .B(_15344_),
    .Y(_15350_));
 sky130_fd_sc_hd__a21oi_2 _37923_ (.A1(_14973_),
    .A2(_14974_),
    .B1(_14967_),
    .Y(_15351_));
 sky130_fd_sc_hd__nand2_2 _37924_ (.A(_15350_),
    .B(_15351_),
    .Y(_15352_));
 sky130_fd_sc_hd__nand3_4 _37925_ (.A(_15339_),
    .B(_15345_),
    .C(_15344_),
    .Y(_15353_));
 sky130_fd_sc_hd__o21ai_1 _37926_ (.A1(_15326_),
    .A2(_15328_),
    .B1(_15329_),
    .Y(_15354_));
 sky130_fd_sc_hd__nand3_2 _37927_ (.A(_15332_),
    .B(_15330_),
    .C(_15327_),
    .Y(_15355_));
 sky130_fd_sc_hd__nand2_2 _37928_ (.A(_15354_),
    .B(_15355_),
    .Y(_15356_));
 sky130_fd_sc_hd__nand3_2 _37929_ (.A(_15352_),
    .B(_15353_),
    .C(_15356_),
    .Y(_15357_));
 sky130_fd_sc_hd__nand3_4 _37930_ (.A(_15323_),
    .B(_15349_),
    .C(_15357_),
    .Y(_15358_));
 sky130_fd_sc_hd__o21a_1 _37931_ (.A1(_15326_),
    .A2(_15328_),
    .B1(_15329_),
    .X(_15359_));
 sky130_vsdinv _37932_ (.A(_15355_),
    .Y(_15360_));
 sky130_fd_sc_hd__o22ai_4 _37933_ (.A1(_15359_),
    .A2(_15360_),
    .B1(_15346_),
    .B2(_15348_),
    .Y(_15361_));
 sky130_fd_sc_hd__o21ai_2 _37934_ (.A1(_14987_),
    .A2(_14977_),
    .B1(_14984_),
    .Y(_15362_));
 sky130_fd_sc_hd__o21ai_1 _37935_ (.A1(_15326_),
    .A2(_15328_),
    .B1(_15330_),
    .Y(_15363_));
 sky130_fd_sc_hd__nand2_2 _37936_ (.A(_15363_),
    .B(_15333_),
    .Y(_15364_));
 sky130_fd_sc_hd__nand3_2 _37937_ (.A(_15352_),
    .B(_15353_),
    .C(_15364_),
    .Y(_15365_));
 sky130_fd_sc_hd__nand3_4 _37938_ (.A(_15361_),
    .B(_15362_),
    .C(_15365_),
    .Y(_15366_));
 sky130_fd_sc_hd__nand2_1 _37939_ (.A(_15358_),
    .B(_15366_),
    .Y(_15367_));
 sky130_fd_sc_hd__o21ai_1 _37940_ (.A1(_14955_),
    .A2(_14956_),
    .B1(_14958_),
    .Y(_15368_));
 sky130_fd_sc_hd__and2_2 _37941_ (.A(_15368_),
    .B(_14959_),
    .X(_15369_));
 sky130_fd_sc_hd__nor2_2 _37942_ (.A(net464),
    .B(_11734_),
    .Y(_15370_));
 sky130_fd_sc_hd__nand2_2 _37943_ (.A(_10383_),
    .B(_07564_),
    .Y(_15371_));
 sky130_fd_sc_hd__a21o_1 _37944_ (.A1(_12818_),
    .A2(_20111_),
    .B1(_15371_),
    .X(_15372_));
 sky130_fd_sc_hd__nand2_1 _37945_ (.A(_10553_),
    .B(_07723_),
    .Y(_15373_));
 sky130_fd_sc_hd__a21o_1 _37946_ (.A1(_11366_),
    .A2(_11062_),
    .B1(_15373_),
    .X(_15374_));
 sky130_fd_sc_hd__nand3b_4 _37947_ (.A_N(_15370_),
    .B(_15372_),
    .C(_15374_),
    .Y(_15375_));
 sky130_fd_sc_hd__nand3b_4 _37948_ (.A_N(_15371_),
    .B(_12818_),
    .C(_20111_),
    .Y(_15376_));
 sky130_fd_sc_hd__nand2_1 _37949_ (.A(_15371_),
    .B(_15373_),
    .Y(_15377_));
 sky130_fd_sc_hd__nand3_4 _37950_ (.A(_15376_),
    .B(_15370_),
    .C(_15377_),
    .Y(_15378_));
 sky130_fd_sc_hd__nand3_4 _37951_ (.A(_15369_),
    .B(_15375_),
    .C(_15378_),
    .Y(_15379_));
 sky130_fd_sc_hd__and2_2 _37952_ (.A(_15007_),
    .B(_15004_),
    .X(_15380_));
 sky130_fd_sc_hd__a21oi_4 _37953_ (.A1(_15375_),
    .A2(_15378_),
    .B1(_15369_),
    .Y(_15381_));
 sky130_fd_sc_hd__nor2_2 _37954_ (.A(_15380_),
    .B(_15381_),
    .Y(_15382_));
 sky130_fd_sc_hd__nand2_1 _37955_ (.A(_15375_),
    .B(_15378_),
    .Y(_15383_));
 sky130_fd_sc_hd__nand2_1 _37956_ (.A(_15368_),
    .B(_14959_),
    .Y(_15384_));
 sky130_fd_sc_hd__nand2_2 _37957_ (.A(_15383_),
    .B(_15384_),
    .Y(_15385_));
 sky130_fd_sc_hd__a21boi_4 _37958_ (.A1(_15385_),
    .A2(_15379_),
    .B1_N(_15380_),
    .Y(_15386_));
 sky130_fd_sc_hd__a21oi_4 _37959_ (.A1(_15379_),
    .A2(_15382_),
    .B1(_15386_),
    .Y(_15387_));
 sky130_fd_sc_hd__nand2_4 _37960_ (.A(_15367_),
    .B(_15387_),
    .Y(_15388_));
 sky130_fd_sc_hd__a21oi_4 _37961_ (.A1(_14980_),
    .A2(_14988_),
    .B1(_14954_),
    .Y(_15389_));
 sky130_fd_sc_hd__a21oi_4 _37962_ (.A1(_14989_),
    .A2(_15018_),
    .B1(_15389_),
    .Y(_15390_));
 sky130_fd_sc_hd__nand2_1 _37963_ (.A(_15385_),
    .B(_15379_),
    .Y(_15391_));
 sky130_fd_sc_hd__nor2_4 _37964_ (.A(_15380_),
    .B(_15391_),
    .Y(_15392_));
 sky130_fd_sc_hd__o211ai_4 _37965_ (.A1(_15386_),
    .A2(_15392_),
    .B1(_15358_),
    .C1(_15366_),
    .Y(_15393_));
 sky130_fd_sc_hd__nand3_4 _37966_ (.A(_15388_),
    .B(_15390_),
    .C(_15393_),
    .Y(_15394_));
 sky130_fd_sc_hd__nand2_1 _37967_ (.A(_14989_),
    .B(_15018_),
    .Y(_15395_));
 sky130_fd_sc_hd__nand2_1 _37968_ (.A(_15395_),
    .B(_14994_),
    .Y(_15396_));
 sky130_fd_sc_hd__o2bb2ai_2 _37969_ (.A1_N(_15358_),
    .A2_N(_15366_),
    .B1(_15386_),
    .B2(_15392_),
    .Y(_15397_));
 sky130_fd_sc_hd__nand3_2 _37970_ (.A(_15387_),
    .B(_15358_),
    .C(_15366_),
    .Y(_15398_));
 sky130_fd_sc_hd__nand3_4 _37971_ (.A(_15396_),
    .B(_15397_),
    .C(_15398_),
    .Y(_15399_));
 sky130_fd_sc_hd__nand2_2 _37972_ (.A(_15008_),
    .B(_15011_),
    .Y(_15400_));
 sky130_fd_sc_hd__a22oi_4 _37973_ (.A1(_13902_),
    .A2(_10716_),
    .B1(_12447_),
    .B2(_10222_),
    .Y(_15401_));
 sky130_fd_sc_hd__and4_4 _37974_ (.A(_12848_),
    .B(_19863_),
    .C(_08881_),
    .D(_09926_),
    .X(_15402_));
 sky130_fd_sc_hd__nand2_4 _37975_ (.A(_07967_),
    .B(_09041_),
    .Y(_15403_));
 sky130_vsdinv _37976_ (.A(_15403_),
    .Y(_15404_));
 sky130_fd_sc_hd__o21ai_2 _37977_ (.A1(_15401_),
    .A2(_15402_),
    .B1(_15404_),
    .Y(_15405_));
 sky130_fd_sc_hd__a21oi_2 _37978_ (.A1(_15037_),
    .A2(_15034_),
    .B1(_15032_),
    .Y(_15406_));
 sky130_fd_sc_hd__nand2_1 _37979_ (.A(_10610_),
    .B(_08450_),
    .Y(_15407_));
 sky130_fd_sc_hd__nand3b_4 _37980_ (.A_N(_15407_),
    .B(_10926_),
    .C(_09044_),
    .Y(_15408_));
 sky130_fd_sc_hd__a22o_2 _37981_ (.A1(_12848_),
    .A2(_08884_),
    .B1(_13497_),
    .B2(_10222_),
    .X(_15409_));
 sky130_fd_sc_hd__nand3_2 _37982_ (.A(_15408_),
    .B(_15409_),
    .C(_15403_),
    .Y(_15410_));
 sky130_fd_sc_hd__nand3_4 _37983_ (.A(_15405_),
    .B(_15406_),
    .C(_15410_),
    .Y(_15411_));
 sky130_fd_sc_hd__o21ai_2 _37984_ (.A1(_15401_),
    .A2(_15402_),
    .B1(_15403_),
    .Y(_15412_));
 sky130_fd_sc_hd__nand3_2 _37985_ (.A(_15408_),
    .B(_15409_),
    .C(_15404_),
    .Y(_15413_));
 sky130_fd_sc_hd__o22ai_4 _37986_ (.A1(_08038_),
    .A2(_15031_),
    .B1(_15033_),
    .B2(_15030_),
    .Y(_15414_));
 sky130_fd_sc_hd__nand3_4 _37987_ (.A(_15412_),
    .B(_15413_),
    .C(_15414_),
    .Y(_15415_));
 sky130_fd_sc_hd__and4_2 _37988_ (.A(_10934_),
    .B(_10944_),
    .C(_20090_),
    .D(_09038_),
    .X(_15416_));
 sky130_fd_sc_hd__nand2_1 _37989_ (.A(_11869_),
    .B(_09899_),
    .Y(_15417_));
 sky130_fd_sc_hd__a22o_1 _37990_ (.A1(_07483_),
    .A2(_10814_),
    .B1(_19874_),
    .B2(_20091_),
    .X(_15418_));
 sky130_fd_sc_hd__nand3b_1 _37991_ (.A_N(_15416_),
    .B(_15417_),
    .C(_15418_),
    .Y(_15419_));
 sky130_fd_sc_hd__a22oi_4 _37992_ (.A1(_07483_),
    .A2(_10814_),
    .B1(_19874_),
    .B2(_09902_),
    .Y(_15420_));
 sky130_vsdinv _37993_ (.A(_15417_),
    .Y(_15421_));
 sky130_fd_sc_hd__o21ai_1 _37994_ (.A1(_15420_),
    .A2(_15416_),
    .B1(_15421_),
    .Y(_15422_));
 sky130_fd_sc_hd__nand2_2 _37995_ (.A(_15419_),
    .B(_15422_),
    .Y(_15423_));
 sky130_fd_sc_hd__a21oi_2 _37996_ (.A1(_15411_),
    .A2(_15415_),
    .B1(_15423_),
    .Y(_15424_));
 sky130_fd_sc_hd__nor3_1 _37997_ (.A(_15421_),
    .B(_15420_),
    .C(_15416_),
    .Y(_15425_));
 sky130_fd_sc_hd__o21a_1 _37998_ (.A1(_15420_),
    .A2(_15416_),
    .B1(_15421_),
    .X(_15426_));
 sky130_fd_sc_hd__o211a_1 _37999_ (.A1(_15425_),
    .A2(_15426_),
    .B1(_15415_),
    .C1(_15411_),
    .X(_15427_));
 sky130_fd_sc_hd__o2bb2ai_4 _38000_ (.A1_N(_15015_),
    .A2_N(_15400_),
    .B1(_15424_),
    .B2(_15427_),
    .Y(_15428_));
 sky130_vsdinv _38001_ (.A(_15415_),
    .Y(_15429_));
 sky130_fd_sc_hd__nand2_2 _38002_ (.A(_15423_),
    .B(_15411_),
    .Y(_15430_));
 sky130_fd_sc_hd__a21oi_4 _38003_ (.A1(_15008_),
    .A2(_15011_),
    .B1(_15012_),
    .Y(_15431_));
 sky130_fd_sc_hd__a21o_1 _38004_ (.A1(_15411_),
    .A2(_15415_),
    .B1(_15423_),
    .X(_15432_));
 sky130_fd_sc_hd__o211ai_4 _38005_ (.A1(_15429_),
    .A2(_15430_),
    .B1(_15431_),
    .C1(_15432_),
    .Y(_15433_));
 sky130_fd_sc_hd__nand2_1 _38006_ (.A(_15054_),
    .B(_15039_),
    .Y(_15434_));
 sky130_fd_sc_hd__nand2_4 _38007_ (.A(_15434_),
    .B(_15043_),
    .Y(_15435_));
 sky130_fd_sc_hd__a21oi_4 _38008_ (.A1(_15428_),
    .A2(_15433_),
    .B1(_15435_),
    .Y(_15436_));
 sky130_fd_sc_hd__nand3_2 _38009_ (.A(_15428_),
    .B(_15433_),
    .C(_15435_),
    .Y(_15437_));
 sky130_vsdinv _38010_ (.A(_15437_),
    .Y(_15438_));
 sky130_fd_sc_hd__o2bb2ai_4 _38011_ (.A1_N(_15394_),
    .A2_N(_15399_),
    .B1(_15436_),
    .B2(_15438_),
    .Y(_15439_));
 sky130_fd_sc_hd__nor2_2 _38012_ (.A(_15436_),
    .B(_15438_),
    .Y(_15440_));
 sky130_fd_sc_hd__nand3_4 _38013_ (.A(_15440_),
    .B(_15399_),
    .C(_15394_),
    .Y(_15441_));
 sky130_fd_sc_hd__nand2_2 _38014_ (.A(_15077_),
    .B(_15027_),
    .Y(_15442_));
 sky130_fd_sc_hd__a21oi_4 _38015_ (.A1(_15439_),
    .A2(_15441_),
    .B1(_15442_),
    .Y(_15443_));
 sky130_fd_sc_hd__nand2_1 _38016_ (.A(_15061_),
    .B(_15066_),
    .Y(_15444_));
 sky130_fd_sc_hd__a31oi_1 _38017_ (.A1(_15020_),
    .A2(_15019_),
    .A3(_15021_),
    .B1(_15444_),
    .Y(_15445_));
 sky130_fd_sc_hd__o211a_2 _38018_ (.A1(_15076_),
    .A2(_15445_),
    .B1(_15441_),
    .C1(_15439_),
    .X(_15446_));
 sky130_fd_sc_hd__o22ai_4 _38019_ (.A1(_15318_),
    .A2(_15320_),
    .B1(_15443_),
    .B2(_15446_),
    .Y(_15447_));
 sky130_fd_sc_hd__a21o_1 _38020_ (.A1(_15439_),
    .A2(_15441_),
    .B1(_15442_),
    .X(_15448_));
 sky130_fd_sc_hd__a21o_1 _38021_ (.A1(_15091_),
    .A2(_15092_),
    .B1(_14812_),
    .X(_15449_));
 sky130_fd_sc_hd__nand3_1 _38022_ (.A(_15091_),
    .B(_14812_),
    .C(_15092_),
    .Y(_15450_));
 sky130_fd_sc_hd__nand2_1 _38023_ (.A(_15449_),
    .B(_15450_),
    .Y(_15451_));
 sky130_fd_sc_hd__nor2_2 _38024_ (.A(_15451_),
    .B(_15116_),
    .Y(_15452_));
 sky130_fd_sc_hd__o2bb2ai_1 _38025_ (.A1_N(_15315_),
    .A2_N(_15311_),
    .B1(_15118_),
    .B2(_15452_),
    .Y(_15453_));
 sky130_fd_sc_hd__nor2_2 _38026_ (.A(_15118_),
    .B(_15452_),
    .Y(_15454_));
 sky130_fd_sc_hd__nand3_1 _38027_ (.A(_15311_),
    .B(_15315_),
    .C(_15454_),
    .Y(_15455_));
 sky130_fd_sc_hd__nand2_2 _38028_ (.A(_15453_),
    .B(_15455_),
    .Y(_15456_));
 sky130_fd_sc_hd__nand3_4 _38029_ (.A(_15442_),
    .B(_15439_),
    .C(_15441_),
    .Y(_15457_));
 sky130_fd_sc_hd__nand3_4 _38030_ (.A(_15448_),
    .B(_15456_),
    .C(_15457_),
    .Y(_15458_));
 sky130_fd_sc_hd__a22oi_4 _38031_ (.A1(_15151_),
    .A2(_15269_),
    .B1(_15447_),
    .B2(_15458_),
    .Y(_15459_));
 sky130_fd_sc_hd__o211a_1 _38032_ (.A1(_15078_),
    .A2(_15141_),
    .B1(_15458_),
    .C1(_15447_),
    .X(_15460_));
 sky130_fd_sc_hd__o22ai_4 _38033_ (.A1(_15267_),
    .A2(_15268_),
    .B1(_15459_),
    .B2(_15460_),
    .Y(_15461_));
 sky130_vsdinv _38034_ (.A(_15072_),
    .Y(_15462_));
 sky130_fd_sc_hd__nand2_1 _38035_ (.A(_15074_),
    .B(_15068_),
    .Y(_15463_));
 sky130_fd_sc_hd__o22ai_4 _38036_ (.A1(_15462_),
    .A2(_15463_),
    .B1(_15135_),
    .B2(_15075_),
    .Y(_15464_));
 sky130_fd_sc_hd__a21o_1 _38037_ (.A1(_15447_),
    .A2(_15458_),
    .B1(_15464_),
    .X(_15465_));
 sky130_fd_sc_hd__nor2_2 _38038_ (.A(_15267_),
    .B(_15268_),
    .Y(_15466_));
 sky130_fd_sc_hd__nand3_4 _38039_ (.A(_15447_),
    .B(_15464_),
    .C(_15458_),
    .Y(_15467_));
 sky130_fd_sc_hd__nand3_4 _38040_ (.A(_15465_),
    .B(_15466_),
    .C(_15467_),
    .Y(_15468_));
 sky130_fd_sc_hd__nand2_1 _38041_ (.A(_15192_),
    .B(_15153_),
    .Y(_15469_));
 sky130_fd_sc_hd__nand2_4 _38042_ (.A(_15469_),
    .B(_15146_),
    .Y(_15470_));
 sky130_fd_sc_hd__a21oi_4 _38043_ (.A1(_15461_),
    .A2(_15468_),
    .B1(_15470_),
    .Y(_15471_));
 sky130_fd_sc_hd__nand2_1 _38044_ (.A(_15466_),
    .B(_15467_),
    .Y(_15472_));
 sky130_fd_sc_hd__o211a_1 _38045_ (.A1(_15459_),
    .A2(_15472_),
    .B1(_15461_),
    .C1(_15470_),
    .X(_15473_));
 sky130_fd_sc_hd__nand2_1 _38046_ (.A(_15195_),
    .B(_15187_),
    .Y(_15474_));
 sky130_fd_sc_hd__nor2_1 _38047_ (.A(_14930_),
    .B(_15474_),
    .Y(_15475_));
 sky130_fd_sc_hd__nand2_2 _38048_ (.A(_15474_),
    .B(_14930_),
    .Y(_15476_));
 sky130_fd_sc_hd__nand2b_4 _38049_ (.A_N(_15475_),
    .B(_15476_),
    .Y(_15477_));
 sky130_fd_sc_hd__o21ai_2 _38050_ (.A1(_15471_),
    .A2(_15473_),
    .B1(_15477_),
    .Y(_15478_));
 sky130_fd_sc_hd__nand2_1 _38051_ (.A(_15198_),
    .B(_15207_),
    .Y(_15479_));
 sky130_fd_sc_hd__nand2_2 _38052_ (.A(_15479_),
    .B(_15202_),
    .Y(_15480_));
 sky130_fd_sc_hd__a21o_1 _38053_ (.A1(_15461_),
    .A2(_15468_),
    .B1(_15470_),
    .X(_15481_));
 sky130_fd_sc_hd__nand3_4 _38054_ (.A(_15470_),
    .B(_15461_),
    .C(_15468_),
    .Y(_15482_));
 sky130_vsdinv _38055_ (.A(_15477_),
    .Y(_15483_));
 sky130_fd_sc_hd__nand3_4 _38056_ (.A(_15481_),
    .B(_15482_),
    .C(_15483_),
    .Y(_15484_));
 sky130_fd_sc_hd__nand3_4 _38057_ (.A(_15478_),
    .B(_15480_),
    .C(_15484_),
    .Y(_15485_));
 sky130_fd_sc_hd__o21ai_4 _38058_ (.A1(_15471_),
    .A2(_15473_),
    .B1(_15483_),
    .Y(_15486_));
 sky130_fd_sc_hd__a21boi_4 _38059_ (.A1(_15198_),
    .A2(_15207_),
    .B1_N(_15202_),
    .Y(_15487_));
 sky130_fd_sc_hd__nand3_4 _38060_ (.A(_15481_),
    .B(_15482_),
    .C(_15477_),
    .Y(_15488_));
 sky130_fd_sc_hd__nand3_4 _38061_ (.A(_15486_),
    .B(_15487_),
    .C(_15488_),
    .Y(_15489_));
 sky130_fd_sc_hd__o2bb2ai_4 _38062_ (.A1_N(_15485_),
    .A2_N(_15489_),
    .B1(_14356_),
    .B2(_15205_),
    .Y(_15490_));
 sky130_fd_sc_hd__nand3_4 _38063_ (.A(_15485_),
    .B(_15489_),
    .C(_15206_),
    .Y(_15491_));
 sky130_fd_sc_hd__a21oi_4 _38064_ (.A1(_15212_),
    .A2(_15213_),
    .B1(_14953_),
    .Y(_15492_));
 sky130_fd_sc_hd__o21ai_4 _38065_ (.A1(_15217_),
    .A2(_15492_),
    .B1(_15214_),
    .Y(_15493_));
 sky130_fd_sc_hd__a21oi_4 _38066_ (.A1(_15490_),
    .A2(_15491_),
    .B1(_15493_),
    .Y(_15494_));
 sky130_fd_sc_hd__nand3_1 _38067_ (.A(_15490_),
    .B(_15493_),
    .C(_15491_),
    .Y(_15495_));
 sky130_vsdinv _38068_ (.A(_15495_),
    .Y(_15496_));
 sky130_fd_sc_hd__nor2_8 _38069_ (.A(_15494_),
    .B(_15496_),
    .Y(_15497_));
 sky130_vsdinv _38070_ (.A(_15219_),
    .Y(_15498_));
 sky130_fd_sc_hd__o21ai_4 _38071_ (.A1(_15498_),
    .A2(_15233_),
    .B1(_15223_),
    .Y(_15499_));
 sky130_fd_sc_hd__xnor2_4 _38072_ (.A(_15497_),
    .B(_15499_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand3_4 _38073_ (.A(_15260_),
    .B(_15265_),
    .C(_15266_),
    .Y(_15500_));
 sky130_fd_sc_hd__nand2_4 _38074_ (.A(_15500_),
    .B(_15265_),
    .Y(_15501_));
 sky130_vsdinv _38075_ (.A(_15501_),
    .Y(_15502_));
 sky130_fd_sc_hd__nor2_8 _38076_ (.A(_13740_),
    .B(_15502_),
    .Y(_15503_));
 sky130_fd_sc_hd__nor2_8 _38077_ (.A(_14930_),
    .B(_15501_),
    .Y(_15504_));
 sky130_fd_sc_hd__nand2_1 _38078_ (.A(_11103_),
    .B(_11587_),
    .Y(_15505_));
 sky130_fd_sc_hd__nand2_1 _38079_ (.A(_19887_),
    .B(_20073_),
    .Y(_15506_));
 sky130_fd_sc_hd__or2_4 _38080_ (.A(_15505_),
    .B(_15506_),
    .X(_15507_));
 sky130_fd_sc_hd__nor2_2 _38081_ (.A(net443),
    .B(_11176_),
    .Y(_15508_));
 sky130_fd_sc_hd__nand2_1 _38082_ (.A(_15505_),
    .B(_15506_),
    .Y(_15509_));
 sky130_fd_sc_hd__nand3_4 _38083_ (.A(_15507_),
    .B(_15508_),
    .C(_15509_),
    .Y(_15510_));
 sky130_fd_sc_hd__a21o_1 _38084_ (.A1(_19888_),
    .A2(_11174_),
    .B1(_15505_),
    .X(_15511_));
 sky130_fd_sc_hd__a21o_1 _38085_ (.A1(_19882_),
    .A2(_10768_),
    .B1(_15506_),
    .X(_15512_));
 sky130_fd_sc_hd__nand3b_4 _38086_ (.A_N(_15508_),
    .B(_15511_),
    .C(_15512_),
    .Y(_15513_));
 sky130_fd_sc_hd__a21o_2 _38087_ (.A1(_15418_),
    .A2(_15421_),
    .B1(_15416_),
    .X(_15514_));
 sky130_fd_sc_hd__a21oi_2 _38088_ (.A1(_15510_),
    .A2(_15513_),
    .B1(_15514_),
    .Y(_15515_));
 sky130_fd_sc_hd__nor2_1 _38089_ (.A(_15417_),
    .B(_15420_),
    .Y(_15516_));
 sky130_fd_sc_hd__o211a_1 _38090_ (.A1(_15416_),
    .A2(_15516_),
    .B1(_15513_),
    .C1(_15510_),
    .X(_15517_));
 sky130_fd_sc_hd__and2_1 _38091_ (.A(_15278_),
    .B(_15276_),
    .X(_15518_));
 sky130_fd_sc_hd__o21ai_4 _38092_ (.A1(_15515_),
    .A2(_15517_),
    .B1(_15518_),
    .Y(_15519_));
 sky130_fd_sc_hd__a21o_2 _38093_ (.A1(_15510_),
    .A2(_15513_),
    .B1(_15514_),
    .X(_15520_));
 sky130_fd_sc_hd__nand2_2 _38094_ (.A(_15278_),
    .B(_15276_),
    .Y(_15521_));
 sky130_fd_sc_hd__nand3_4 _38095_ (.A(_15510_),
    .B(_15514_),
    .C(_15513_),
    .Y(_15522_));
 sky130_fd_sc_hd__nand3_4 _38096_ (.A(_15520_),
    .B(_15521_),
    .C(_15522_),
    .Y(_15523_));
 sky130_fd_sc_hd__o21ai_4 _38097_ (.A1(_15284_),
    .A2(_15280_),
    .B1(_15287_),
    .Y(_15524_));
 sky130_fd_sc_hd__a21oi_4 _38098_ (.A1(_15519_),
    .A2(_15523_),
    .B1(_15524_),
    .Y(_15525_));
 sky130_fd_sc_hd__nand2_1 _38099_ (.A(_15520_),
    .B(_15521_),
    .Y(_15526_));
 sky130_fd_sc_hd__o211a_1 _38100_ (.A1(_15517_),
    .A2(_15526_),
    .B1(_15524_),
    .C1(_15519_),
    .X(_15527_));
 sky130_fd_sc_hd__and3_2 _38101_ (.A(_14806_),
    .B(_19893_),
    .C(_06359_),
    .X(_15528_));
 sky130_fd_sc_hd__o21ai_4 _38102_ (.A1(_19894_),
    .A2(_19897_),
    .B1(_18687_),
    .Y(_15529_));
 sky130_fd_sc_hd__o21ai_2 _38103_ (.A1(_13271_),
    .A2(_15297_),
    .B1(_15294_),
    .Y(_15530_));
 sky130_fd_sc_hd__o21bai_4 _38104_ (.A1(_15528_),
    .A2(_15529_),
    .B1_N(_15530_),
    .Y(_15531_));
 sky130_vsdinv _38105_ (.A(_15528_),
    .Y(_15532_));
 sky130_fd_sc_hd__nand3b_4 _38106_ (.A_N(_15529_),
    .B(_15530_),
    .C(_15532_),
    .Y(_15533_));
 sky130_fd_sc_hd__nand2_1 _38107_ (.A(_15531_),
    .B(_15533_),
    .Y(_15534_));
 sky130_fd_sc_hd__nand2_1 _38108_ (.A(_15534_),
    .B(_14812_),
    .Y(_15535_));
 sky130_fd_sc_hd__nand3_1 _38109_ (.A(_15531_),
    .B(_14844_),
    .C(_15533_),
    .Y(_15536_));
 sky130_fd_sc_hd__and2_1 _38110_ (.A(_15535_),
    .B(_15536_),
    .X(_15537_));
 sky130_fd_sc_hd__o21ai_2 _38111_ (.A1(_15525_),
    .A2(_15527_),
    .B1(_15537_),
    .Y(_15538_));
 sky130_fd_sc_hd__a21boi_2 _38112_ (.A1(_15428_),
    .A2(_15435_),
    .B1_N(_15433_),
    .Y(_15539_));
 sky130_fd_sc_hd__a21o_1 _38113_ (.A1(_15519_),
    .A2(_15523_),
    .B1(_15524_),
    .X(_15540_));
 sky130_fd_sc_hd__nand3_4 _38114_ (.A(_15519_),
    .B(_15524_),
    .C(_15523_),
    .Y(_15541_));
 sky130_fd_sc_hd__nand2_1 _38115_ (.A(_15535_),
    .B(_15536_),
    .Y(_15542_));
 sky130_fd_sc_hd__nand3_2 _38116_ (.A(_15540_),
    .B(_15541_),
    .C(_15542_),
    .Y(_15543_));
 sky130_fd_sc_hd__nand3_4 _38117_ (.A(_15538_),
    .B(_15539_),
    .C(_15543_),
    .Y(_15544_));
 sky130_fd_sc_hd__o21ai_2 _38118_ (.A1(_15525_),
    .A2(_15527_),
    .B1(_15542_),
    .Y(_15545_));
 sky130_fd_sc_hd__nand2_1 _38119_ (.A(_15437_),
    .B(_15433_),
    .Y(_15546_));
 sky130_fd_sc_hd__nand3_2 _38120_ (.A(_15537_),
    .B(_15540_),
    .C(_15541_),
    .Y(_15547_));
 sky130_fd_sc_hd__nand3_4 _38121_ (.A(_15545_),
    .B(_15546_),
    .C(_15547_),
    .Y(_15548_));
 sky130_fd_sc_hd__nor2_2 _38122_ (.A(_15305_),
    .B(_15290_),
    .Y(_15549_));
 sky130_fd_sc_hd__or2_4 _38123_ (.A(_15291_),
    .B(_15549_),
    .X(_15550_));
 sky130_fd_sc_hd__a21oi_4 _38124_ (.A1(_15544_),
    .A2(_15548_),
    .B1(_15550_),
    .Y(_15551_));
 sky130_fd_sc_hd__nand3_4 _38125_ (.A(_15550_),
    .B(_15544_),
    .C(_15548_),
    .Y(_15552_));
 sky130_vsdinv _38126_ (.A(_15552_),
    .Y(_15553_));
 sky130_fd_sc_hd__nand2_1 _38127_ (.A(_15387_),
    .B(_15358_),
    .Y(_15554_));
 sky130_fd_sc_hd__nand2_2 _38128_ (.A(_15554_),
    .B(_15366_),
    .Y(_15555_));
 sky130_fd_sc_hd__nor2_1 _38129_ (.A(_09321_),
    .B(_11057_),
    .Y(_15556_));
 sky130_vsdinv _38130_ (.A(_15556_),
    .Y(_15557_));
 sky130_fd_sc_hd__nand2_2 _38131_ (.A(_11794_),
    .B(_06976_),
    .Y(_15558_));
 sky130_fd_sc_hd__nand2_2 _38132_ (.A(_19840_),
    .B(_20118_),
    .Y(_15559_));
 sky130_fd_sc_hd__nor2_2 _38133_ (.A(_15558_),
    .B(_15559_),
    .Y(_15560_));
 sky130_fd_sc_hd__nand2_2 _38134_ (.A(_15558_),
    .B(_15559_),
    .Y(_15561_));
 sky130_vsdinv _38135_ (.A(_15561_),
    .Y(_15562_));
 sky130_fd_sc_hd__nor2_1 _38136_ (.A(_15560_),
    .B(_15562_),
    .Y(_15563_));
 sky130_fd_sc_hd__nor2_2 _38137_ (.A(_15557_),
    .B(_15563_),
    .Y(_15564_));
 sky130_fd_sc_hd__and2_1 _38138_ (.A(_15563_),
    .B(_15557_),
    .X(_15565_));
 sky130_fd_sc_hd__nand3_4 _38139_ (.A(_10973_),
    .B(_11783_),
    .C(_06714_),
    .Y(_15566_));
 sky130_fd_sc_hd__nor2_4 _38140_ (.A(_10941_),
    .B(_15566_),
    .Y(_15567_));
 sky130_fd_sc_hd__a22oi_4 _38141_ (.A1(_13138_),
    .A2(_11093_),
    .B1(_06440_),
    .B2(_13139_),
    .Y(_15568_));
 sky130_fd_sc_hd__nand2_4 _38142_ (.A(_10573_),
    .B(_20126_),
    .Y(_15569_));
 sky130_fd_sc_hd__o21ai_4 _38143_ (.A1(_15567_),
    .A2(_15568_),
    .B1(_15569_),
    .Y(_15570_));
 sky130_vsdinv _38144_ (.A(_15569_),
    .Y(_15571_));
 sky130_fd_sc_hd__o2bb2ai_4 _38145_ (.A1_N(_13138_),
    .A2_N(_12846_),
    .B1(_10941_),
    .B2(_13142_),
    .Y(_15572_));
 sky130_fd_sc_hd__o211ai_4 _38146_ (.A1(_20134_),
    .A2(_15566_),
    .B1(_15571_),
    .C1(_15572_),
    .Y(_15573_));
 sky130_fd_sc_hd__o21ai_4 _38147_ (.A1(_15338_),
    .A2(_15337_),
    .B1(_15341_),
    .Y(_15574_));
 sky130_fd_sc_hd__a21oi_4 _38148_ (.A1(_15570_),
    .A2(_15573_),
    .B1(_15574_),
    .Y(_15575_));
 sky130_fd_sc_hd__a21oi_4 _38149_ (.A1(_15342_),
    .A2(_15343_),
    .B1(_15336_),
    .Y(_15576_));
 sky130_fd_sc_hd__nand2_2 _38150_ (.A(_15570_),
    .B(_15573_),
    .Y(_15577_));
 sky130_fd_sc_hd__nor2_4 _38151_ (.A(_15576_),
    .B(_15577_),
    .Y(_15578_));
 sky130_fd_sc_hd__o22ai_4 _38152_ (.A1(_15564_),
    .A2(_15565_),
    .B1(_15575_),
    .B2(_15578_),
    .Y(_15579_));
 sky130_vsdinv _38153_ (.A(_15344_),
    .Y(_15580_));
 sky130_fd_sc_hd__nand2_1 _38154_ (.A(_15339_),
    .B(_15345_),
    .Y(_15581_));
 sky130_fd_sc_hd__a2bb2oi_4 _38155_ (.A1_N(_15580_),
    .A2_N(_15581_),
    .B1(_15364_),
    .B2(_15352_),
    .Y(_15582_));
 sky130_fd_sc_hd__nand2_2 _38156_ (.A(_15577_),
    .B(_15576_),
    .Y(_15583_));
 sky130_fd_sc_hd__nand3_4 _38157_ (.A(_15570_),
    .B(_15574_),
    .C(_15573_),
    .Y(_15584_));
 sky130_fd_sc_hd__o21ai_2 _38158_ (.A1(_15560_),
    .A2(_15562_),
    .B1(_15557_),
    .Y(_15585_));
 sky130_fd_sc_hd__nand3b_2 _38159_ (.A_N(_15560_),
    .B(_15556_),
    .C(_15561_),
    .Y(_15586_));
 sky130_fd_sc_hd__nand2_4 _38160_ (.A(_15585_),
    .B(_15586_),
    .Y(_15587_));
 sky130_fd_sc_hd__nand3_4 _38161_ (.A(_15583_),
    .B(_15584_),
    .C(_15587_),
    .Y(_15588_));
 sky130_fd_sc_hd__nand3_4 _38162_ (.A(_15579_),
    .B(_15582_),
    .C(_15588_),
    .Y(_15589_));
 sky130_fd_sc_hd__o21ai_2 _38163_ (.A1(_15575_),
    .A2(_15578_),
    .B1(_15587_),
    .Y(_15590_));
 sky130_fd_sc_hd__o21ai_2 _38164_ (.A1(_15356_),
    .A2(_15346_),
    .B1(_15353_),
    .Y(_15591_));
 sky130_fd_sc_hd__nand3b_2 _38165_ (.A_N(_15587_),
    .B(_15583_),
    .C(_15584_),
    .Y(_15592_));
 sky130_fd_sc_hd__nand3_4 _38166_ (.A(_15590_),
    .B(_15591_),
    .C(_15592_),
    .Y(_15593_));
 sky130_fd_sc_hd__buf_2 _38167_ (.A(_19851_),
    .X(_15594_));
 sky130_fd_sc_hd__nand2_1 _38168_ (.A(_19848_),
    .B(_10711_),
    .Y(_15595_));
 sky130_fd_sc_hd__a21o_1 _38169_ (.A1(_15594_),
    .A2(_13758_),
    .B1(_15595_),
    .X(_15596_));
 sky130_fd_sc_hd__buf_2 _38170_ (.A(_11826_),
    .X(_15597_));
 sky130_fd_sc_hd__nand2_2 _38171_ (.A(_11371_),
    .B(_10343_),
    .Y(_15598_));
 sky130_fd_sc_hd__a21o_1 _38172_ (.A1(_15597_),
    .A2(_11492_),
    .B1(_15598_),
    .X(_15599_));
 sky130_fd_sc_hd__nand2_1 _38173_ (.A(_19855_),
    .B(_11085_),
    .Y(_15600_));
 sky130_fd_sc_hd__nand3_4 _38174_ (.A(_15596_),
    .B(_15599_),
    .C(_15600_),
    .Y(_15601_));
 sky130_fd_sc_hd__nand3_2 _38175_ (.A(_15597_),
    .B(_15594_),
    .C(_11492_),
    .Y(_15602_));
 sky130_fd_sc_hd__nand2_1 _38176_ (.A(_15595_),
    .B(_15598_),
    .Y(_15603_));
 sky130_fd_sc_hd__o2111ai_4 _38177_ (.A1(_09733_),
    .A2(_15602_),
    .B1(_19855_),
    .C1(_11085_),
    .D1(_15603_),
    .Y(_15604_));
 sky130_fd_sc_hd__nand2_1 _38178_ (.A(_15601_),
    .B(_15604_),
    .Y(_15605_));
 sky130_fd_sc_hd__o21ai_1 _38179_ (.A1(_15324_),
    .A2(_15325_),
    .B1(_15329_),
    .Y(_15606_));
 sky130_fd_sc_hd__nand2_2 _38180_ (.A(_15606_),
    .B(_15327_),
    .Y(_15607_));
 sky130_fd_sc_hd__nand2_4 _38181_ (.A(_15605_),
    .B(_15607_),
    .Y(_15608_));
 sky130_fd_sc_hd__nand3b_4 _38182_ (.A_N(_15607_),
    .B(_15601_),
    .C(_15604_),
    .Y(_15609_));
 sky130_fd_sc_hd__nand2_4 _38183_ (.A(_15378_),
    .B(_15376_),
    .Y(_15610_));
 sky130_fd_sc_hd__a21oi_4 _38184_ (.A1(_15608_),
    .A2(_15609_),
    .B1(_15610_),
    .Y(_15611_));
 sky130_fd_sc_hd__nand3_2 _38185_ (.A(_15608_),
    .B(_15609_),
    .C(_15610_),
    .Y(_15612_));
 sky130_vsdinv _38186_ (.A(_15612_),
    .Y(_15613_));
 sky130_fd_sc_hd__o2bb2ai_4 _38187_ (.A1_N(_15589_),
    .A2_N(_15593_),
    .B1(_15611_),
    .B2(_15613_),
    .Y(_15614_));
 sky130_fd_sc_hd__and2_1 _38188_ (.A(_15378_),
    .B(_15376_),
    .X(_15615_));
 sky130_fd_sc_hd__a21boi_4 _38189_ (.A1(_15601_),
    .A2(_15604_),
    .B1_N(_15607_),
    .Y(_15616_));
 sky130_fd_sc_hd__nor2_4 _38190_ (.A(_15615_),
    .B(_15616_),
    .Y(_15617_));
 sky130_fd_sc_hd__a21oi_4 _38191_ (.A1(_15617_),
    .A2(_15609_),
    .B1(_15611_),
    .Y(_15618_));
 sky130_fd_sc_hd__nand3_4 _38192_ (.A(_15593_),
    .B(_15589_),
    .C(_15618_),
    .Y(_15619_));
 sky130_fd_sc_hd__nand3_4 _38193_ (.A(_15555_),
    .B(_15614_),
    .C(_15619_),
    .Y(_15620_));
 sky130_fd_sc_hd__a21oi_1 _38194_ (.A1(_15324_),
    .A2(_15325_),
    .B1(_15329_),
    .Y(_15621_));
 sky130_fd_sc_hd__o211a_2 _38195_ (.A1(_15326_),
    .A2(_15621_),
    .B1(_15604_),
    .C1(_15601_),
    .X(_15622_));
 sky130_fd_sc_hd__o21ai_1 _38196_ (.A1(_15616_),
    .A2(_15622_),
    .B1(_15615_),
    .Y(_15623_));
 sky130_fd_sc_hd__nand2_2 _38197_ (.A(_15623_),
    .B(_15612_),
    .Y(_15624_));
 sky130_fd_sc_hd__a21o_1 _38198_ (.A1(_15593_),
    .A2(_15589_),
    .B1(_15624_),
    .X(_15625_));
 sky130_fd_sc_hd__a21boi_4 _38199_ (.A1(_15387_),
    .A2(_15358_),
    .B1_N(_15366_),
    .Y(_15626_));
 sky130_fd_sc_hd__nand3_2 _38200_ (.A(_15593_),
    .B(_15589_),
    .C(_15624_),
    .Y(_15627_));
 sky130_fd_sc_hd__nand3_4 _38201_ (.A(_15625_),
    .B(_15626_),
    .C(_15627_),
    .Y(_15628_));
 sky130_vsdinv _38202_ (.A(_15411_),
    .Y(_15629_));
 sky130_fd_sc_hd__nor2_2 _38203_ (.A(_15423_),
    .B(_15429_),
    .Y(_15630_));
 sky130_fd_sc_hd__nand2_1 _38204_ (.A(_15408_),
    .B(_15403_),
    .Y(_15631_));
 sky130_fd_sc_hd__nand2_4 _38205_ (.A(_10433_),
    .B(_08446_),
    .Y(_15632_));
 sky130_fd_sc_hd__nand2_4 _38206_ (.A(_10620_),
    .B(_09041_),
    .Y(_15633_));
 sky130_fd_sc_hd__nor2_4 _38207_ (.A(_15632_),
    .B(_15633_),
    .Y(_15634_));
 sky130_fd_sc_hd__nor2_4 _38208_ (.A(_07822_),
    .B(_11549_),
    .Y(_15635_));
 sky130_fd_sc_hd__nand2_4 _38209_ (.A(_15632_),
    .B(_15633_),
    .Y(_15636_));
 sky130_fd_sc_hd__nand3b_4 _38210_ (.A_N(_15634_),
    .B(_15635_),
    .C(_15636_),
    .Y(_15637_));
 sky130_fd_sc_hd__a21o_1 _38211_ (.A1(_10926_),
    .A2(_09493_),
    .B1(_15632_),
    .X(_15638_));
 sky130_fd_sc_hd__a21o_1 _38212_ (.A1(_10917_),
    .A2(_10811_),
    .B1(_15633_),
    .X(_15639_));
 sky130_fd_sc_hd__o211ai_4 _38213_ (.A1(_07822_),
    .A2(_11557_),
    .B1(_15638_),
    .C1(_15639_),
    .Y(_15640_));
 sky130_fd_sc_hd__a22oi_4 _38214_ (.A1(_15631_),
    .A2(_15409_),
    .B1(_15637_),
    .B2(_15640_),
    .Y(_15641_));
 sky130_fd_sc_hd__nor2_4 _38215_ (.A(_15403_),
    .B(_15401_),
    .Y(_15642_));
 sky130_fd_sc_hd__o211a_2 _38216_ (.A1(_15402_),
    .A2(_15642_),
    .B1(_15640_),
    .C1(_15637_),
    .X(_15643_));
 sky130_fd_sc_hd__nand2_1 _38217_ (.A(_12864_),
    .B(_11210_),
    .Y(_15644_));
 sky130_fd_sc_hd__nand2_1 _38218_ (.A(_07902_),
    .B(_09899_),
    .Y(_15645_));
 sky130_fd_sc_hd__nor2_1 _38219_ (.A(_15644_),
    .B(_15645_),
    .Y(_15646_));
 sky130_fd_sc_hd__nor2_1 _38220_ (.A(_07141_),
    .B(_09775_),
    .Y(_15647_));
 sky130_vsdinv _38221_ (.A(_15647_),
    .Y(_15648_));
 sky130_fd_sc_hd__nand2_1 _38222_ (.A(_15644_),
    .B(_15645_),
    .Y(_15649_));
 sky130_fd_sc_hd__nand3b_1 _38223_ (.A_N(_15646_),
    .B(_15648_),
    .C(_15649_),
    .Y(_15650_));
 sky130_vsdinv _38224_ (.A(_15649_),
    .Y(_15651_));
 sky130_fd_sc_hd__o21ai_1 _38225_ (.A1(_15646_),
    .A2(_15651_),
    .B1(_15647_),
    .Y(_15652_));
 sky130_fd_sc_hd__nand2_2 _38226_ (.A(_15650_),
    .B(_15652_),
    .Y(_15653_));
 sky130_fd_sc_hd__o21bai_4 _38227_ (.A1(_15641_),
    .A2(_15643_),
    .B1_N(_15653_),
    .Y(_15654_));
 sky130_fd_sc_hd__nand2_1 _38228_ (.A(_15637_),
    .B(_15640_),
    .Y(_15655_));
 sky130_fd_sc_hd__nor2_1 _38229_ (.A(_15402_),
    .B(_15642_),
    .Y(_15656_));
 sky130_fd_sc_hd__nand2_2 _38230_ (.A(_15655_),
    .B(_15656_),
    .Y(_15657_));
 sky130_fd_sc_hd__o211ai_4 _38231_ (.A1(_15402_),
    .A2(_15642_),
    .B1(_15640_),
    .C1(_15637_),
    .Y(_15658_));
 sky130_fd_sc_hd__nand3_4 _38232_ (.A(_15657_),
    .B(_15658_),
    .C(_15653_),
    .Y(_15659_));
 sky130_fd_sc_hd__o21ai_4 _38233_ (.A1(_15380_),
    .A2(_15381_),
    .B1(_15379_),
    .Y(_15660_));
 sky130_fd_sc_hd__a21oi_4 _38234_ (.A1(_15654_),
    .A2(_15659_),
    .B1(_15660_),
    .Y(_15661_));
 sky130_fd_sc_hd__nand2_1 _38235_ (.A(_15657_),
    .B(_15653_),
    .Y(_15662_));
 sky130_fd_sc_hd__o211a_2 _38236_ (.A1(_15643_),
    .A2(_15662_),
    .B1(_15660_),
    .C1(_15654_),
    .X(_15663_));
 sky130_fd_sc_hd__o22ai_4 _38237_ (.A1(_15629_),
    .A2(_15630_),
    .B1(_15661_),
    .B2(_15663_),
    .Y(_15664_));
 sky130_vsdinv _38238_ (.A(_15664_),
    .Y(_15665_));
 sky130_fd_sc_hd__a21o_1 _38239_ (.A1(_15654_),
    .A2(_15659_),
    .B1(_15660_),
    .X(_15666_));
 sky130_fd_sc_hd__nand3_2 _38240_ (.A(_15654_),
    .B(_15660_),
    .C(_15659_),
    .Y(_15667_));
 sky130_fd_sc_hd__nand2_2 _38241_ (.A(_15430_),
    .B(_15415_),
    .Y(_15668_));
 sky130_fd_sc_hd__nand3_2 _38242_ (.A(_15666_),
    .B(_15667_),
    .C(_15668_),
    .Y(_15669_));
 sky130_vsdinv _38243_ (.A(_15669_),
    .Y(_15670_));
 sky130_fd_sc_hd__o2bb2ai_4 _38244_ (.A1_N(_15620_),
    .A2_N(_15628_),
    .B1(_15665_),
    .B2(_15670_),
    .Y(_15671_));
 sky130_fd_sc_hd__nand2_1 _38245_ (.A(_15666_),
    .B(_15668_),
    .Y(_15672_));
 sky130_fd_sc_hd__o21a_1 _38246_ (.A1(_15663_),
    .A2(_15672_),
    .B1(_15664_),
    .X(_15673_));
 sky130_fd_sc_hd__nand3_4 _38247_ (.A(_15673_),
    .B(_15628_),
    .C(_15620_),
    .Y(_15674_));
 sky130_fd_sc_hd__nand2_1 _38248_ (.A(_15440_),
    .B(_15394_),
    .Y(_15675_));
 sky130_fd_sc_hd__nand2_2 _38249_ (.A(_15675_),
    .B(_15399_),
    .Y(_15676_));
 sky130_fd_sc_hd__a21oi_4 _38250_ (.A1(_15671_),
    .A2(_15674_),
    .B1(_15676_),
    .Y(_15677_));
 sky130_vsdinv _38251_ (.A(_15399_),
    .Y(_15678_));
 sky130_fd_sc_hd__a21o_1 _38252_ (.A1(_15428_),
    .A2(_15433_),
    .B1(_15435_),
    .X(_15679_));
 sky130_fd_sc_hd__nand2_1 _38253_ (.A(_15679_),
    .B(_15437_),
    .Y(_15680_));
 sky130_fd_sc_hd__a31oi_4 _38254_ (.A1(_15390_),
    .A2(_15388_),
    .A3(_15393_),
    .B1(_15680_),
    .Y(_15681_));
 sky130_fd_sc_hd__o211a_2 _38255_ (.A1(_15678_),
    .A2(_15681_),
    .B1(_15674_),
    .C1(_15671_),
    .X(_15682_));
 sky130_fd_sc_hd__o22ai_4 _38256_ (.A1(_15551_),
    .A2(_15553_),
    .B1(_15677_),
    .B2(_15682_),
    .Y(_15683_));
 sky130_fd_sc_hd__o2bb2ai_1 _38257_ (.A1_N(_15315_),
    .A2_N(_15311_),
    .B1(_15116_),
    .B2(_15316_),
    .Y(_15684_));
 sky130_fd_sc_hd__nand2_1 _38258_ (.A(_15684_),
    .B(_15319_),
    .Y(_15685_));
 sky130_fd_sc_hd__o21ai_4 _38259_ (.A1(_15443_),
    .A2(_15685_),
    .B1(_15457_),
    .Y(_15686_));
 sky130_fd_sc_hd__nand2_1 _38260_ (.A(_15671_),
    .B(_15674_),
    .Y(_15687_));
 sky130_fd_sc_hd__nor2_2 _38261_ (.A(_15678_),
    .B(_15681_),
    .Y(_15688_));
 sky130_fd_sc_hd__nand2_2 _38262_ (.A(_15687_),
    .B(_15688_),
    .Y(_15689_));
 sky130_fd_sc_hd__o21a_1 _38263_ (.A1(_15291_),
    .A2(_15549_),
    .B1(_15544_),
    .X(_15690_));
 sky130_fd_sc_hd__a21oi_4 _38264_ (.A1(_15690_),
    .A2(_15548_),
    .B1(_15551_),
    .Y(_15691_));
 sky130_fd_sc_hd__nand3_4 _38265_ (.A(_15676_),
    .B(_15671_),
    .C(_15674_),
    .Y(_15692_));
 sky130_fd_sc_hd__nand3_4 _38266_ (.A(_15689_),
    .B(_15691_),
    .C(_15692_),
    .Y(_15693_));
 sky130_fd_sc_hd__nand3_4 _38267_ (.A(_15683_),
    .B(_15686_),
    .C(_15693_),
    .Y(_15694_));
 sky130_fd_sc_hd__o21ai_2 _38268_ (.A1(_15677_),
    .A2(_15682_),
    .B1(_15691_),
    .Y(_15695_));
 sky130_fd_sc_hd__a21oi_4 _38269_ (.A1(_15448_),
    .A2(_15456_),
    .B1(_15446_),
    .Y(_15696_));
 sky130_fd_sc_hd__nand2_1 _38270_ (.A(_15544_),
    .B(_15548_),
    .Y(_15697_));
 sky130_fd_sc_hd__nor2_1 _38271_ (.A(_15291_),
    .B(_15549_),
    .Y(_15698_));
 sky130_fd_sc_hd__nand2_1 _38272_ (.A(_15697_),
    .B(_15698_),
    .Y(_15699_));
 sky130_fd_sc_hd__nand2_2 _38273_ (.A(_15699_),
    .B(_15552_),
    .Y(_15700_));
 sky130_fd_sc_hd__nand3_2 _38274_ (.A(_15689_),
    .B(_15700_),
    .C(_15692_),
    .Y(_15701_));
 sky130_fd_sc_hd__nand3_4 _38275_ (.A(_15695_),
    .B(_15696_),
    .C(_15701_),
    .Y(_15702_));
 sky130_vsdinv _38276_ (.A(_15262_),
    .Y(_15703_));
 sky130_fd_sc_hd__nand3_4 _38277_ (.A(_15165_),
    .B(_15300_),
    .C(_15303_),
    .Y(_15704_));
 sky130_fd_sc_hd__nand2_1 _38278_ (.A(_15303_),
    .B(_15300_),
    .Y(_15705_));
 sky130_fd_sc_hd__nand3_4 _38279_ (.A(_15705_),
    .B(_15164_),
    .C(_15163_),
    .Y(_15706_));
 sky130_fd_sc_hd__a21o_1 _38280_ (.A1(_15704_),
    .A2(_15706_),
    .B1(_15244_),
    .X(_15707_));
 sky130_fd_sc_hd__nand3_4 _38281_ (.A(_15704_),
    .B(_15244_),
    .C(_15706_),
    .Y(_15708_));
 sky130_fd_sc_hd__nand2_2 _38282_ (.A(_15707_),
    .B(_15708_),
    .Y(_15709_));
 sky130_fd_sc_hd__o21a_1 _38283_ (.A1(_15165_),
    .A2(_15238_),
    .B1(_15252_),
    .X(_15710_));
 sky130_fd_sc_hd__nand2_1 _38284_ (.A(_15709_),
    .B(_15710_),
    .Y(_15711_));
 sky130_fd_sc_hd__nand2_2 _38285_ (.A(_15252_),
    .B(_15241_),
    .Y(_15712_));
 sky130_fd_sc_hd__nand3_4 _38286_ (.A(_15712_),
    .B(_15707_),
    .C(_15708_),
    .Y(_15713_));
 sky130_fd_sc_hd__nand2_1 _38287_ (.A(_15711_),
    .B(_15713_),
    .Y(_15714_));
 sky130_fd_sc_hd__nand2_1 _38288_ (.A(_15714_),
    .B(_14009_),
    .Y(_15715_));
 sky130_fd_sc_hd__nand2_1 _38289_ (.A(_15308_),
    .B(_15309_),
    .Y(_15716_));
 sky130_fd_sc_hd__a21oi_2 _38290_ (.A1(_15716_),
    .A2(_15305_),
    .B1(_15313_),
    .Y(_15717_));
 sky130_fd_sc_hd__a22oi_4 _38291_ (.A1(_15717_),
    .A2(_15310_),
    .B1(_15315_),
    .B2(_15317_),
    .Y(_15718_));
 sky130_fd_sc_hd__nand3_2 _38292_ (.A(_15711_),
    .B(_14303_),
    .C(_15713_),
    .Y(_15719_));
 sky130_fd_sc_hd__nand3_4 _38293_ (.A(_15715_),
    .B(_15718_),
    .C(_15719_),
    .Y(_15720_));
 sky130_fd_sc_hd__and3_1 _38294_ (.A(_15306_),
    .B(_15307_),
    .C(_15310_),
    .X(_15721_));
 sky130_fd_sc_hd__a31oi_4 _38295_ (.A1(_15312_),
    .A2(_15313_),
    .A3(_15314_),
    .B1(_15454_),
    .Y(_15722_));
 sky130_fd_sc_hd__a21oi_4 _38296_ (.A1(_15709_),
    .A2(_15710_),
    .B1(_14303_),
    .Y(_15723_));
 sky130_fd_sc_hd__nand2_1 _38297_ (.A(_15723_),
    .B(_15713_),
    .Y(_15724_));
 sky130_fd_sc_hd__nand2_1 _38298_ (.A(_15714_),
    .B(_13679_),
    .Y(_15725_));
 sky130_fd_sc_hd__o211ai_4 _38299_ (.A1(_15721_),
    .A2(_15722_),
    .B1(_15724_),
    .C1(_15725_),
    .Y(_15726_));
 sky130_fd_sc_hd__o211a_1 _38300_ (.A1(_15261_),
    .A2(_15703_),
    .B1(_15720_),
    .C1(_15726_),
    .X(_15727_));
 sky130_fd_sc_hd__nand2_2 _38301_ (.A(_15262_),
    .B(_15256_),
    .Y(_15728_));
 sky130_fd_sc_hd__a21oi_2 _38302_ (.A1(_15726_),
    .A2(_15720_),
    .B1(_15728_),
    .Y(_15729_));
 sky130_fd_sc_hd__o2bb2ai_2 _38303_ (.A1_N(_15694_),
    .A2_N(_15702_),
    .B1(_15727_),
    .B2(_15729_),
    .Y(_15730_));
 sky130_vsdinv _38304_ (.A(_15458_),
    .Y(_15731_));
 sky130_fd_sc_hd__nand2_1 _38305_ (.A(_15447_),
    .B(_15464_),
    .Y(_15732_));
 sky130_fd_sc_hd__nand2_1 _38306_ (.A(_15260_),
    .B(_15265_),
    .Y(_15733_));
 sky130_vsdinv _38307_ (.A(_15266_),
    .Y(_15734_));
 sky130_fd_sc_hd__nand2_1 _38308_ (.A(_15733_),
    .B(_15734_),
    .Y(_15735_));
 sky130_fd_sc_hd__nand2_1 _38309_ (.A(_15735_),
    .B(_15500_),
    .Y(_15736_));
 sky130_fd_sc_hd__o22ai_4 _38310_ (.A1(_15731_),
    .A2(_15732_),
    .B1(_15736_),
    .B2(_15459_),
    .Y(_15737_));
 sky130_fd_sc_hd__nor2_2 _38311_ (.A(_15729_),
    .B(_15727_),
    .Y(_15738_));
 sky130_fd_sc_hd__nand3_2 _38312_ (.A(_15738_),
    .B(_15694_),
    .C(_15702_),
    .Y(_15739_));
 sky130_fd_sc_hd__nand3_4 _38313_ (.A(_15730_),
    .B(_15737_),
    .C(_15739_),
    .Y(_15740_));
 sky130_fd_sc_hd__nand2_1 _38314_ (.A(_15702_),
    .B(_15694_),
    .Y(_15741_));
 sky130_fd_sc_hd__nand2_1 _38315_ (.A(_15741_),
    .B(_15738_),
    .Y(_15742_));
 sky130_fd_sc_hd__o21ai_1 _38316_ (.A1(_15267_),
    .A2(_15268_),
    .B1(_15467_),
    .Y(_15743_));
 sky130_fd_sc_hd__nand2_1 _38317_ (.A(_15743_),
    .B(_15465_),
    .Y(_15744_));
 sky130_fd_sc_hd__nand2_1 _38318_ (.A(_15726_),
    .B(_15720_),
    .Y(_15745_));
 sky130_vsdinv _38319_ (.A(_15728_),
    .Y(_15746_));
 sky130_fd_sc_hd__nand2_1 _38320_ (.A(_15745_),
    .B(_15746_),
    .Y(_15747_));
 sky130_fd_sc_hd__nand3_1 _38321_ (.A(_15726_),
    .B(_15720_),
    .C(_15728_),
    .Y(_15748_));
 sky130_fd_sc_hd__nand2_2 _38322_ (.A(_15747_),
    .B(_15748_),
    .Y(_15749_));
 sky130_fd_sc_hd__nand3_2 _38323_ (.A(_15749_),
    .B(_15702_),
    .C(_15694_),
    .Y(_15750_));
 sky130_fd_sc_hd__nand3_4 _38324_ (.A(_15742_),
    .B(_15744_),
    .C(_15750_),
    .Y(_15751_));
 sky130_fd_sc_hd__o211ai_4 _38325_ (.A1(_15503_),
    .A2(_15504_),
    .B1(_15740_),
    .C1(_15751_),
    .Y(_15752_));
 sky130_fd_sc_hd__nor2_1 _38326_ (.A(_14931_),
    .B(_15502_),
    .Y(_15753_));
 sky130_fd_sc_hd__buf_6 _38327_ (.A(_13740_),
    .X(_15754_));
 sky130_fd_sc_hd__nor2_1 _38328_ (.A(_15754_),
    .B(_15501_),
    .Y(_15755_));
 sky130_fd_sc_hd__o2bb2ai_2 _38329_ (.A1_N(_15740_),
    .A2_N(_15751_),
    .B1(_15753_),
    .B2(_15755_),
    .Y(_15756_));
 sky130_fd_sc_hd__o2111ai_4 _38330_ (.A1(_15477_),
    .A2(_15471_),
    .B1(_15482_),
    .C1(_15752_),
    .D1(_15756_),
    .Y(_15757_));
 sky130_vsdinv _38331_ (.A(_15468_),
    .Y(_15758_));
 sky130_fd_sc_hd__nand2_1 _38332_ (.A(_15470_),
    .B(_15461_),
    .Y(_15759_));
 sky130_fd_sc_hd__o22ai_4 _38333_ (.A1(_15758_),
    .A2(_15759_),
    .B1(_15477_),
    .B2(_15471_),
    .Y(_15760_));
 sky130_fd_sc_hd__o2bb2ai_2 _38334_ (.A1_N(_15740_),
    .A2_N(_15751_),
    .B1(_15503_),
    .B2(_15504_),
    .Y(_15761_));
 sky130_fd_sc_hd__nor2_4 _38335_ (.A(_15504_),
    .B(_15503_),
    .Y(_15762_));
 sky130_fd_sc_hd__nand3_4 _38336_ (.A(_15751_),
    .B(_15740_),
    .C(_15762_),
    .Y(_15763_));
 sky130_fd_sc_hd__nand3_4 _38337_ (.A(_15760_),
    .B(_15761_),
    .C(_15763_),
    .Y(_15764_));
 sky130_vsdinv _38338_ (.A(_15476_),
    .Y(_15765_));
 sky130_fd_sc_hd__a21oi_1 _38339_ (.A1(_15757_),
    .A2(_15764_),
    .B1(_15765_),
    .Y(_15766_));
 sky130_fd_sc_hd__and3_1 _38340_ (.A(_15757_),
    .B(_15764_),
    .C(_15765_),
    .X(_15767_));
 sky130_vsdinv _38341_ (.A(_15206_),
    .Y(_15768_));
 sky130_fd_sc_hd__a31oi_4 _38342_ (.A1(_15486_),
    .A2(_15487_),
    .A3(_15488_),
    .B1(_15768_),
    .Y(_15769_));
 sky130_fd_sc_hd__and3_1 _38343_ (.A(_15478_),
    .B(_15480_),
    .C(_15484_),
    .X(_15770_));
 sky130_fd_sc_hd__nor2_1 _38344_ (.A(_15769_),
    .B(_15770_),
    .Y(_15771_));
 sky130_fd_sc_hd__o21ai_2 _38345_ (.A1(_15766_),
    .A2(_15767_),
    .B1(_15771_),
    .Y(_15772_));
 sky130_fd_sc_hd__nand3_2 _38346_ (.A(_15757_),
    .B(_15764_),
    .C(_15765_),
    .Y(_15773_));
 sky130_fd_sc_hd__a21o_1 _38347_ (.A1(_15757_),
    .A2(_15764_),
    .B1(_15765_),
    .X(_15774_));
 sky130_fd_sc_hd__o211ai_4 _38348_ (.A1(_15769_),
    .A2(_15770_),
    .B1(_15773_),
    .C1(_15774_),
    .Y(_15775_));
 sky130_fd_sc_hd__nand2_2 _38349_ (.A(_15772_),
    .B(_15775_),
    .Y(_15776_));
 sky130_vsdinv _38350_ (.A(_15491_),
    .Y(_15777_));
 sky130_fd_sc_hd__nand2_1 _38351_ (.A(_15490_),
    .B(_15493_),
    .Y(_15778_));
 sky130_fd_sc_hd__a21o_1 _38352_ (.A1(_15490_),
    .A2(_15491_),
    .B1(_15493_),
    .X(_15779_));
 sky130_fd_sc_hd__o2111ai_4 _38353_ (.A1(_15777_),
    .A2(_15778_),
    .B1(_15223_),
    .C1(_15219_),
    .D1(_15779_),
    .Y(_15780_));
 sky130_vsdinv _38354_ (.A(_15780_),
    .Y(_15781_));
 sky130_fd_sc_hd__a21o_1 _38355_ (.A1(_15219_),
    .A2(_15495_),
    .B1(_15494_),
    .X(_15782_));
 sky130_fd_sc_hd__a21boi_4 _38356_ (.A1(_15233_),
    .A2(_15781_),
    .B1_N(_15782_),
    .Y(_15783_));
 sky130_fd_sc_hd__xor2_4 _38357_ (.A(_15776_),
    .B(_15783_),
    .X(_02665_));
 sky130_vsdinv _38358_ (.A(_15713_),
    .Y(_15784_));
 sky130_fd_sc_hd__nor2_4 _38359_ (.A(_15784_),
    .B(_15723_),
    .Y(_15785_));
 sky130_fd_sc_hd__nand2_1 _38360_ (.A(_15552_),
    .B(_15548_),
    .Y(_15786_));
 sky130_fd_sc_hd__nor2_8 _38361_ (.A(_13271_),
    .B(_15532_),
    .Y(_15787_));
 sky130_fd_sc_hd__a21oi_4 _38362_ (.A1(_15531_),
    .A2(_15533_),
    .B1(_14844_),
    .Y(_15788_));
 sky130_fd_sc_hd__nor2_2 _38363_ (.A(_15162_),
    .B(_15160_),
    .Y(_15789_));
 sky130_fd_sc_hd__nor2_4 _38364_ (.A(_14279_),
    .B(_15158_),
    .Y(_15790_));
 sky130_fd_sc_hd__nor2_1 _38365_ (.A(_15789_),
    .B(_15790_),
    .Y(_15791_));
 sky130_fd_sc_hd__o21bai_1 _38366_ (.A1(_15787_),
    .A2(_15788_),
    .B1_N(_15791_),
    .Y(_15792_));
 sky130_vsdinv _38367_ (.A(_15787_),
    .Y(_15793_));
 sky130_fd_sc_hd__nand3_1 _38368_ (.A(_15535_),
    .B(_15793_),
    .C(_15791_),
    .Y(_15794_));
 sky130_fd_sc_hd__nand2_1 _38369_ (.A(_15792_),
    .B(_15794_),
    .Y(_15795_));
 sky130_fd_sc_hd__nand3b_4 _38370_ (.A_N(_15795_),
    .B(_15706_),
    .C(_15708_),
    .Y(_15796_));
 sky130_fd_sc_hd__nand2_1 _38371_ (.A(_15708_),
    .B(_15706_),
    .Y(_15797_));
 sky130_fd_sc_hd__nand2_2 _38372_ (.A(_15797_),
    .B(_15795_),
    .Y(_15798_));
 sky130_fd_sc_hd__a21o_1 _38373_ (.A1(_15796_),
    .A2(_15798_),
    .B1(_14310_),
    .X(_15799_));
 sky130_fd_sc_hd__nand3_4 _38374_ (.A(_15796_),
    .B(_15798_),
    .C(_14310_),
    .Y(_15800_));
 sky130_fd_sc_hd__nand3_4 _38375_ (.A(_15786_),
    .B(_15799_),
    .C(_15800_),
    .Y(_15801_));
 sky130_fd_sc_hd__nand2_2 _38376_ (.A(_15799_),
    .B(_15800_),
    .Y(_15802_));
 sky130_fd_sc_hd__a21boi_4 _38377_ (.A1(_15550_),
    .A2(_15544_),
    .B1_N(_15548_),
    .Y(_15803_));
 sky130_fd_sc_hd__nand2_4 _38378_ (.A(_15802_),
    .B(_15803_),
    .Y(_15804_));
 sky130_fd_sc_hd__nand2_1 _38379_ (.A(_15801_),
    .B(_15804_),
    .Y(_15805_));
 sky130_fd_sc_hd__nor2_4 _38380_ (.A(_15785_),
    .B(_15805_),
    .Y(_15806_));
 sky130_vsdinv _38381_ (.A(_15785_),
    .Y(_15807_));
 sky130_fd_sc_hd__a21oi_4 _38382_ (.A1(_15801_),
    .A2(_15804_),
    .B1(_15807_),
    .Y(_15808_));
 sky130_fd_sc_hd__nand2_2 _38383_ (.A(_11103_),
    .B(_20073_),
    .Y(_15809_));
 sky130_fd_sc_hd__nand2_2 _38384_ (.A(_11094_),
    .B(_20069_),
    .Y(_15810_));
 sky130_fd_sc_hd__nor2_1 _38385_ (.A(_15809_),
    .B(_15810_),
    .Y(_15811_));
 sky130_fd_sc_hd__and2_1 _38386_ (.A(_15809_),
    .B(_15810_),
    .X(_15812_));
 sky130_fd_sc_hd__nand2_4 _38387_ (.A(_18686_),
    .B(net456),
    .Y(_15813_));
 sky130_fd_sc_hd__o21ai_2 _38388_ (.A1(_15811_),
    .A2(_15812_),
    .B1(_15813_),
    .Y(_15814_));
 sky130_fd_sc_hd__or2_2 _38389_ (.A(_15809_),
    .B(_15810_),
    .X(_15815_));
 sky130_vsdinv _38390_ (.A(_15813_),
    .Y(_15816_));
 sky130_fd_sc_hd__nand2_1 _38391_ (.A(_15809_),
    .B(_15810_),
    .Y(_15817_));
 sky130_fd_sc_hd__nand3_4 _38392_ (.A(_15815_),
    .B(_15816_),
    .C(_15817_),
    .Y(_15818_));
 sky130_fd_sc_hd__a31o_2 _38393_ (.A1(_15649_),
    .A2(_19879_),
    .A3(_20083_),
    .B1(_15646_),
    .X(_15819_));
 sky130_fd_sc_hd__a21o_2 _38394_ (.A1(_15814_),
    .A2(_15818_),
    .B1(_15819_),
    .X(_15820_));
 sky130_fd_sc_hd__nand3_4 _38395_ (.A(_15814_),
    .B(_15818_),
    .C(_15819_),
    .Y(_15821_));
 sky130_fd_sc_hd__nand2_4 _38396_ (.A(_15510_),
    .B(_15507_),
    .Y(_15822_));
 sky130_fd_sc_hd__a21oi_4 _38397_ (.A1(_15820_),
    .A2(_15821_),
    .B1(_15822_),
    .Y(_15823_));
 sky130_fd_sc_hd__nand3_4 _38398_ (.A(_15820_),
    .B(_15821_),
    .C(_15822_),
    .Y(_15824_));
 sky130_fd_sc_hd__nand2_2 _38399_ (.A(_15518_),
    .B(_15522_),
    .Y(_15825_));
 sky130_fd_sc_hd__nand3_4 _38400_ (.A(_15824_),
    .B(_15520_),
    .C(_15825_),
    .Y(_15826_));
 sky130_fd_sc_hd__nor2_8 _38401_ (.A(_15823_),
    .B(_15826_),
    .Y(_15827_));
 sky130_fd_sc_hd__a21o_2 _38402_ (.A1(_15820_),
    .A2(_15821_),
    .B1(_15822_),
    .X(_15828_));
 sky130_fd_sc_hd__nand2_1 _38403_ (.A(_15825_),
    .B(_15520_),
    .Y(_15829_));
 sky130_fd_sc_hd__a21boi_4 _38404_ (.A1(_15828_),
    .A2(_15824_),
    .B1_N(_15829_),
    .Y(_15830_));
 sky130_fd_sc_hd__a21o_2 _38405_ (.A1(_15082_),
    .A2(_15529_),
    .B1(_15787_),
    .X(_15831_));
 sky130_fd_sc_hd__nor2_8 _38406_ (.A(_14844_),
    .B(_15831_),
    .Y(_15832_));
 sky130_fd_sc_hd__and2_4 _38407_ (.A(_15831_),
    .B(_14844_),
    .X(_15833_));
 sky130_fd_sc_hd__nor2_8 _38408_ (.A(_15832_),
    .B(_15833_),
    .Y(_15834_));
 sky130_fd_sc_hd__clkbuf_4 _38409_ (.A(_15834_),
    .X(_15835_));
 sky130_fd_sc_hd__o21ai_2 _38410_ (.A1(_15827_),
    .A2(_15830_),
    .B1(_15835_),
    .Y(_15836_));
 sky130_fd_sc_hd__a21oi_4 _38411_ (.A1(_15666_),
    .A2(_15668_),
    .B1(_15663_),
    .Y(_15837_));
 sky130_fd_sc_hd__nand2_1 _38412_ (.A(_15828_),
    .B(_15824_),
    .Y(_15838_));
 sky130_fd_sc_hd__nand2_2 _38413_ (.A(_15838_),
    .B(_15829_),
    .Y(_15839_));
 sky130_fd_sc_hd__or2_4 _38414_ (.A(_15832_),
    .B(_15833_),
    .X(_15840_));
 sky130_fd_sc_hd__nand3b_4 _38415_ (.A_N(_15829_),
    .B(_15828_),
    .C(_15824_),
    .Y(_15841_));
 sky130_fd_sc_hd__nand3_4 _38416_ (.A(_15839_),
    .B(_15840_),
    .C(_15841_),
    .Y(_15842_));
 sky130_fd_sc_hd__nand3_4 _38417_ (.A(_15836_),
    .B(_15837_),
    .C(_15842_),
    .Y(_15843_));
 sky130_fd_sc_hd__o22ai_4 _38418_ (.A1(_15833_),
    .A2(_15832_),
    .B1(_15827_),
    .B2(_15830_),
    .Y(_15844_));
 sky130_fd_sc_hd__nand3_2 _38419_ (.A(_15839_),
    .B(_15835_),
    .C(_15841_),
    .Y(_15845_));
 sky130_vsdinv _38420_ (.A(_15668_),
    .Y(_15846_));
 sky130_fd_sc_hd__o21ai_2 _38421_ (.A1(_15846_),
    .A2(_15661_),
    .B1(_15667_),
    .Y(_15847_));
 sky130_fd_sc_hd__nand3_4 _38422_ (.A(_15844_),
    .B(_15845_),
    .C(_15847_),
    .Y(_15848_));
 sky130_fd_sc_hd__nand2_1 _38423_ (.A(_15537_),
    .B(_15540_),
    .Y(_15849_));
 sky130_fd_sc_hd__nand2_2 _38424_ (.A(_15849_),
    .B(_15541_),
    .Y(_15850_));
 sky130_fd_sc_hd__and3_1 _38425_ (.A(_15843_),
    .B(_15848_),
    .C(_15850_),
    .X(_15851_));
 sky130_fd_sc_hd__a21oi_4 _38426_ (.A1(_15843_),
    .A2(_15848_),
    .B1(_15850_),
    .Y(_15852_));
 sky130_vsdinv _38427_ (.A(_15662_),
    .Y(_15853_));
 sky130_fd_sc_hd__nand2_1 _38428_ (.A(_11396_),
    .B(_12304_),
    .Y(_15854_));
 sky130_fd_sc_hd__a21o_2 _38429_ (.A1(_19864_),
    .A2(_13451_),
    .B1(_15854_),
    .X(_15855_));
 sky130_fd_sc_hd__nand2_1 _38430_ (.A(_12855_),
    .B(_13451_),
    .Y(_15856_));
 sky130_fd_sc_hd__a21o_2 _38431_ (.A1(_19860_),
    .A2(_12304_),
    .B1(_15856_),
    .X(_15857_));
 sky130_fd_sc_hd__nand2_4 _38432_ (.A(_19867_),
    .B(_20092_),
    .Y(_15858_));
 sky130_fd_sc_hd__a21o_1 _38433_ (.A1(_15855_),
    .A2(_15857_),
    .B1(_15858_),
    .X(_15859_));
 sky130_fd_sc_hd__nand3_4 _38434_ (.A(_15855_),
    .B(_15857_),
    .C(_15858_),
    .Y(_15860_));
 sky130_fd_sc_hd__a31o_2 _38435_ (.A1(_15636_),
    .A2(_19868_),
    .A3(_20095_),
    .B1(_15634_),
    .X(_15861_));
 sky130_fd_sc_hd__a21oi_4 _38436_ (.A1(_15859_),
    .A2(_15860_),
    .B1(_15861_),
    .Y(_15862_));
 sky130_fd_sc_hd__a21oi_4 _38437_ (.A1(_15635_),
    .A2(_15636_),
    .B1(_15634_),
    .Y(_15863_));
 sky130_fd_sc_hd__a21oi_4 _38438_ (.A1(_15855_),
    .A2(_15857_),
    .B1(_15858_),
    .Y(_15864_));
 sky130_fd_sc_hd__and3_1 _38439_ (.A(_15855_),
    .B(_15857_),
    .C(_15858_),
    .X(_15865_));
 sky130_fd_sc_hd__nor3_4 _38440_ (.A(_15863_),
    .B(_15864_),
    .C(_15865_),
    .Y(_15866_));
 sky130_fd_sc_hd__nand2_4 _38441_ (.A(_12298_),
    .B(_10262_),
    .Y(_15867_));
 sky130_fd_sc_hd__a22o_1 _38442_ (.A1(_10935_),
    .A2(_11934_),
    .B1(_10936_),
    .B2(_12298_),
    .X(_15868_));
 sky130_fd_sc_hd__nor2_4 _38443_ (.A(_07141_),
    .B(_12688_),
    .Y(_15869_));
 sky130_fd_sc_hd__o211a_1 _38444_ (.A1(_12219_),
    .A2(_15867_),
    .B1(_15868_),
    .C1(_15869_),
    .X(_15870_));
 sky130_fd_sc_hd__buf_2 _38445_ (.A(_12219_),
    .X(_15871_));
 sky130_fd_sc_hd__o21ai_4 _38446_ (.A1(_15871_),
    .A2(_15867_),
    .B1(_15868_),
    .Y(_15872_));
 sky130_fd_sc_hd__o21a_1 _38447_ (.A1(_07141_),
    .A2(_11181_),
    .B1(_15872_),
    .X(_15873_));
 sky130_fd_sc_hd__nor2_4 _38448_ (.A(_15870_),
    .B(_15873_),
    .Y(_15874_));
 sky130_fd_sc_hd__o21ai_2 _38449_ (.A1(_15862_),
    .A2(_15866_),
    .B1(_15874_),
    .Y(_15875_));
 sky130_fd_sc_hd__a21oi_4 _38450_ (.A1(_15608_),
    .A2(_15610_),
    .B1(_15622_),
    .Y(_15876_));
 sky130_fd_sc_hd__o21ai_2 _38451_ (.A1(_15864_),
    .A2(_15865_),
    .B1(_15863_),
    .Y(_15877_));
 sky130_fd_sc_hd__xor2_4 _38452_ (.A(_15869_),
    .B(_15872_),
    .X(_15878_));
 sky130_fd_sc_hd__nand3_4 _38453_ (.A(_15859_),
    .B(_15861_),
    .C(_15860_),
    .Y(_15879_));
 sky130_fd_sc_hd__nand3_2 _38454_ (.A(_15877_),
    .B(_15878_),
    .C(_15879_),
    .Y(_15880_));
 sky130_fd_sc_hd__nand3_4 _38455_ (.A(_15875_),
    .B(_15876_),
    .C(_15880_),
    .Y(_15881_));
 sky130_fd_sc_hd__nand2_4 _38456_ (.A(_15877_),
    .B(_15874_),
    .Y(_15882_));
 sky130_fd_sc_hd__o21ai_2 _38457_ (.A1(_15862_),
    .A2(_15866_),
    .B1(_15878_),
    .Y(_15883_));
 sky130_fd_sc_hd__o221ai_4 _38458_ (.A1(_15622_),
    .A2(_15617_),
    .B1(_15866_),
    .B2(_15882_),
    .C1(_15883_),
    .Y(_15884_));
 sky130_fd_sc_hd__o211a_1 _38459_ (.A1(_15643_),
    .A2(_15853_),
    .B1(_15881_),
    .C1(_15884_),
    .X(_15885_));
 sky130_fd_sc_hd__nand2_2 _38460_ (.A(_15662_),
    .B(_15658_),
    .Y(_15886_));
 sky130_fd_sc_hd__a21oi_4 _38461_ (.A1(_15884_),
    .A2(_15881_),
    .B1(_15886_),
    .Y(_15887_));
 sky130_fd_sc_hd__nand2_2 _38462_ (.A(_19855_),
    .B(_20103_),
    .Y(_15888_));
 sky130_fd_sc_hd__nand2_1 _38463_ (.A(_15597_),
    .B(_20108_),
    .Y(_15889_));
 sky130_fd_sc_hd__nand2_1 _38464_ (.A(_15594_),
    .B(_20105_),
    .Y(_15890_));
 sky130_fd_sc_hd__or2_2 _38465_ (.A(_15889_),
    .B(_15890_),
    .X(_15891_));
 sky130_fd_sc_hd__nand2_1 _38466_ (.A(_15889_),
    .B(_15890_),
    .Y(_15892_));
 sky130_fd_sc_hd__nand3b_4 _38467_ (.A_N(_15888_),
    .B(_15891_),
    .C(_15892_),
    .Y(_15893_));
 sky130_fd_sc_hd__nor2_2 _38468_ (.A(_15889_),
    .B(_15890_),
    .Y(_15894_));
 sky130_fd_sc_hd__and2_1 _38469_ (.A(_15889_),
    .B(_15890_),
    .X(_15895_));
 sky130_fd_sc_hd__o21ai_4 _38470_ (.A1(_15894_),
    .A2(_15895_),
    .B1(_15888_),
    .Y(_15896_));
 sky130_fd_sc_hd__clkbuf_4 _38471_ (.A(_19844_),
    .X(_15897_));
 sky130_fd_sc_hd__a31o_2 _38472_ (.A1(_15561_),
    .A2(_15897_),
    .A3(_20116_),
    .B1(_15560_),
    .X(_15898_));
 sky130_fd_sc_hd__a21o_1 _38473_ (.A1(_15893_),
    .A2(_15896_),
    .B1(_15898_),
    .X(_15899_));
 sky130_fd_sc_hd__nand3_4 _38474_ (.A(_15893_),
    .B(_15896_),
    .C(_15898_),
    .Y(_15900_));
 sky130_fd_sc_hd__o21a_1 _38475_ (.A1(_15595_),
    .A2(_15598_),
    .B1(_15604_),
    .X(_15901_));
 sky130_vsdinv _38476_ (.A(_15901_),
    .Y(_15902_));
 sky130_fd_sc_hd__a21oi_2 _38477_ (.A1(_15899_),
    .A2(_15900_),
    .B1(_15902_),
    .Y(_15903_));
 sky130_fd_sc_hd__and3_1 _38478_ (.A(_15899_),
    .B(_15902_),
    .C(_15900_),
    .X(_15904_));
 sky130_fd_sc_hd__nand3_4 _38479_ (.A(_13837_),
    .B(_13138_),
    .C(_20127_),
    .Y(_15905_));
 sky130_fd_sc_hd__nor2_4 _38480_ (.A(_20131_),
    .B(_15905_),
    .Y(_15906_));
 sky130_fd_sc_hd__buf_2 _38481_ (.A(_13138_),
    .X(_15907_));
 sky130_fd_sc_hd__buf_2 _38482_ (.A(_13837_),
    .X(_15908_));
 sky130_fd_sc_hd__a22oi_4 _38483_ (.A1(_15907_),
    .A2(_20127_),
    .B1(_07995_),
    .B2(_15908_),
    .Y(_15909_));
 sky130_fd_sc_hd__nand2_2 _38484_ (.A(_19833_),
    .B(_20124_),
    .Y(_15910_));
 sky130_fd_sc_hd__o21ai_2 _38485_ (.A1(_15906_),
    .A2(_15909_),
    .B1(_15910_),
    .Y(_15911_));
 sky130_fd_sc_hd__o21bai_4 _38486_ (.A1(_15569_),
    .A2(_15568_),
    .B1_N(_15567_),
    .Y(_15912_));
 sky130_vsdinv _38487_ (.A(_15910_),
    .Y(_15913_));
 sky130_fd_sc_hd__buf_2 _38488_ (.A(_11275_),
    .X(_15914_));
 sky130_vsdinv _38489_ (.A(_10575_),
    .Y(_15915_));
 sky130_fd_sc_hd__buf_2 _38490_ (.A(_15915_),
    .X(_15916_));
 sky130_fd_sc_hd__o22ai_4 _38491_ (.A1(_20131_),
    .A2(_15914_),
    .B1(_15916_),
    .B2(_11096_),
    .Y(_15917_));
 sky130_fd_sc_hd__o211ai_4 _38492_ (.A1(_20131_),
    .A2(_15905_),
    .B1(_15913_),
    .C1(_15917_),
    .Y(_15918_));
 sky130_fd_sc_hd__nand3_4 _38493_ (.A(_15911_),
    .B(_15912_),
    .C(_15918_),
    .Y(_15919_));
 sky130_fd_sc_hd__o21ai_2 _38494_ (.A1(_15906_),
    .A2(_15909_),
    .B1(_15913_),
    .Y(_15920_));
 sky130_fd_sc_hd__nand3b_2 _38495_ (.A_N(_15906_),
    .B(_15910_),
    .C(_15917_),
    .Y(_15921_));
 sky130_fd_sc_hd__a21oi_4 _38496_ (.A1(_15572_),
    .A2(_15571_),
    .B1(_15567_),
    .Y(_15922_));
 sky130_fd_sc_hd__nand3_4 _38497_ (.A(_15920_),
    .B(_15921_),
    .C(_15922_),
    .Y(_15923_));
 sky130_fd_sc_hd__buf_2 _38498_ (.A(_09997_),
    .X(_15924_));
 sky130_fd_sc_hd__buf_2 _38499_ (.A(_19841_),
    .X(_15925_));
 sky130_fd_sc_hd__a22oi_4 _38500_ (.A1(_15924_),
    .A2(_20120_),
    .B1(_15925_),
    .B2(_20115_),
    .Y(_15926_));
 sky130_fd_sc_hd__and4_1 _38501_ (.A(_19836_),
    .B(_19841_),
    .C(_20115_),
    .D(_20119_),
    .X(_15927_));
 sky130_fd_sc_hd__nor2_2 _38502_ (.A(_15926_),
    .B(_15927_),
    .Y(_15928_));
 sky130_fd_sc_hd__buf_4 _38503_ (.A(_10340_),
    .X(_15929_));
 sky130_fd_sc_hd__nor2_2 _38504_ (.A(_09321_),
    .B(_15929_),
    .Y(_15930_));
 sky130_fd_sc_hd__and2_1 _38505_ (.A(_15928_),
    .B(_15930_),
    .X(_15931_));
 sky130_fd_sc_hd__nor2_2 _38506_ (.A(_15930_),
    .B(_15928_),
    .Y(_15932_));
 sky130_fd_sc_hd__o2bb2ai_4 _38507_ (.A1_N(_15919_),
    .A2_N(_15923_),
    .B1(_15931_),
    .B2(_15932_),
    .Y(_15933_));
 sky130_fd_sc_hd__o21ai_1 _38508_ (.A1(_09321_),
    .A2(_15929_),
    .B1(_15928_),
    .Y(_15934_));
 sky130_fd_sc_hd__o21ai_1 _38509_ (.A1(_15926_),
    .A2(_15927_),
    .B1(_15930_),
    .Y(_15935_));
 sky130_fd_sc_hd__nand2_2 _38510_ (.A(_15934_),
    .B(_15935_),
    .Y(_15936_));
 sky130_fd_sc_hd__nand3_4 _38511_ (.A(_15936_),
    .B(_15923_),
    .C(_15919_),
    .Y(_15937_));
 sky130_vsdinv _38512_ (.A(_15573_),
    .Y(_15938_));
 sky130_fd_sc_hd__nand2_1 _38513_ (.A(_15570_),
    .B(_15574_),
    .Y(_15939_));
 sky130_fd_sc_hd__o22ai_4 _38514_ (.A1(_15938_),
    .A2(_15939_),
    .B1(_15587_),
    .B2(_15575_),
    .Y(_15940_));
 sky130_fd_sc_hd__a21oi_2 _38515_ (.A1(_15933_),
    .A2(_15937_),
    .B1(_15940_),
    .Y(_15941_));
 sky130_fd_sc_hd__and3_1 _38516_ (.A(_15911_),
    .B(_15912_),
    .C(_15918_),
    .X(_15942_));
 sky130_fd_sc_hd__nand2_2 _38517_ (.A(_15936_),
    .B(_15923_),
    .Y(_15943_));
 sky130_fd_sc_hd__o211a_4 _38518_ (.A1(_15942_),
    .A2(_15943_),
    .B1(_15933_),
    .C1(_15940_),
    .X(_15944_));
 sky130_fd_sc_hd__o22ai_4 _38519_ (.A1(_15903_),
    .A2(_15904_),
    .B1(_15941_),
    .B2(_15944_),
    .Y(_15945_));
 sky130_fd_sc_hd__a21o_1 _38520_ (.A1(_15933_),
    .A2(_15937_),
    .B1(_15940_),
    .X(_15946_));
 sky130_fd_sc_hd__a21oi_4 _38521_ (.A1(_15893_),
    .A2(_15896_),
    .B1(_15898_),
    .Y(_15947_));
 sky130_fd_sc_hd__and3_1 _38522_ (.A(_15893_),
    .B(_15896_),
    .C(_15898_),
    .X(_15948_));
 sky130_fd_sc_hd__o21ai_1 _38523_ (.A1(_15947_),
    .A2(_15948_),
    .B1(_15902_),
    .Y(_15949_));
 sky130_fd_sc_hd__nand3_1 _38524_ (.A(_15899_),
    .B(_15901_),
    .C(_15900_),
    .Y(_15950_));
 sky130_fd_sc_hd__nand2_2 _38525_ (.A(_15949_),
    .B(_15950_),
    .Y(_15951_));
 sky130_fd_sc_hd__nand3_2 _38526_ (.A(_15940_),
    .B(_15933_),
    .C(_15937_),
    .Y(_15952_));
 sky130_fd_sc_hd__nand3_4 _38527_ (.A(_15946_),
    .B(_15951_),
    .C(_15952_),
    .Y(_15953_));
 sky130_fd_sc_hd__nand2_1 _38528_ (.A(_15589_),
    .B(_15618_),
    .Y(_15954_));
 sky130_fd_sc_hd__nand2_2 _38529_ (.A(_15954_),
    .B(_15593_),
    .Y(_15955_));
 sky130_fd_sc_hd__a21oi_4 _38530_ (.A1(_15945_),
    .A2(_15953_),
    .B1(_15955_),
    .Y(_15956_));
 sky130_fd_sc_hd__a21oi_1 _38531_ (.A1(_15579_),
    .A2(_15588_),
    .B1(_15582_),
    .Y(_15957_));
 sky130_fd_sc_hd__a31oi_1 _38532_ (.A1(_15579_),
    .A2(_15582_),
    .A3(_15588_),
    .B1(_15624_),
    .Y(_15958_));
 sky130_fd_sc_hd__o211a_1 _38533_ (.A1(_15957_),
    .A2(_15958_),
    .B1(_15953_),
    .C1(_15945_),
    .X(_15959_));
 sky130_fd_sc_hd__o22ai_4 _38534_ (.A1(_15885_),
    .A2(_15887_),
    .B1(_15956_),
    .B2(_15959_),
    .Y(_15960_));
 sky130_fd_sc_hd__a21o_1 _38535_ (.A1(_15945_),
    .A2(_15953_),
    .B1(_15955_),
    .X(_15961_));
 sky130_fd_sc_hd__nor2_2 _38536_ (.A(_15887_),
    .B(_15885_),
    .Y(_15962_));
 sky130_fd_sc_hd__nand3_4 _38537_ (.A(_15955_),
    .B(_15945_),
    .C(_15953_),
    .Y(_15963_));
 sky130_fd_sc_hd__nand3_4 _38538_ (.A(_15961_),
    .B(_15962_),
    .C(_15963_),
    .Y(_15964_));
 sky130_fd_sc_hd__nand2_2 _38539_ (.A(_15664_),
    .B(_15669_),
    .Y(_15965_));
 sky130_fd_sc_hd__a21oi_4 _38540_ (.A1(_15614_),
    .A2(_15619_),
    .B1(_15555_),
    .Y(_15966_));
 sky130_fd_sc_hd__o21ai_4 _38541_ (.A1(_15965_),
    .A2(_15966_),
    .B1(_15620_),
    .Y(_15967_));
 sky130_fd_sc_hd__a21oi_2 _38542_ (.A1(_15960_),
    .A2(_15964_),
    .B1(_15967_),
    .Y(_15968_));
 sky130_fd_sc_hd__nand2_1 _38543_ (.A(_15614_),
    .B(_15619_),
    .Y(_15969_));
 sky130_fd_sc_hd__nor2_1 _38544_ (.A(_15626_),
    .B(_15969_),
    .Y(_15970_));
 sky130_fd_sc_hd__a21oi_1 _38545_ (.A1(_15969_),
    .A2(_15626_),
    .B1(_15965_),
    .Y(_15971_));
 sky130_fd_sc_hd__o211a_1 _38546_ (.A1(_15970_),
    .A2(_15971_),
    .B1(_15964_),
    .C1(_15960_),
    .X(_15972_));
 sky130_fd_sc_hd__o22ai_4 _38547_ (.A1(_15851_),
    .A2(_15852_),
    .B1(_15968_),
    .B2(_15972_),
    .Y(_15973_));
 sky130_fd_sc_hd__a21o_1 _38548_ (.A1(_15960_),
    .A2(_15964_),
    .B1(_15967_),
    .X(_15974_));
 sky130_fd_sc_hd__and2_1 _38549_ (.A(_15849_),
    .B(_15541_),
    .X(_15975_));
 sky130_fd_sc_hd__a31oi_2 _38550_ (.A1(_15837_),
    .A2(_15836_),
    .A3(_15842_),
    .B1(_15975_),
    .Y(_15976_));
 sky130_fd_sc_hd__a21oi_2 _38551_ (.A1(_15976_),
    .A2(_15848_),
    .B1(_15852_),
    .Y(_15977_));
 sky130_fd_sc_hd__nand3_4 _38552_ (.A(_15967_),
    .B(_15960_),
    .C(_15964_),
    .Y(_15978_));
 sky130_fd_sc_hd__nand3_4 _38553_ (.A(_15974_),
    .B(_15977_),
    .C(_15978_),
    .Y(_15979_));
 sky130_fd_sc_hd__o21ai_4 _38554_ (.A1(_15700_),
    .A2(_15677_),
    .B1(_15692_),
    .Y(_15980_));
 sky130_fd_sc_hd__a21oi_4 _38555_ (.A1(_15973_),
    .A2(_15979_),
    .B1(_15980_),
    .Y(_15981_));
 sky130_fd_sc_hd__a21oi_1 _38556_ (.A1(_15688_),
    .A2(_15687_),
    .B1(_15700_),
    .Y(_15982_));
 sky130_fd_sc_hd__o211a_1 _38557_ (.A1(_15682_),
    .A2(_15982_),
    .B1(_15979_),
    .C1(_15973_),
    .X(_15983_));
 sky130_fd_sc_hd__o22ai_4 _38558_ (.A1(_15806_),
    .A2(_15808_),
    .B1(_15981_),
    .B2(_15983_),
    .Y(_15984_));
 sky130_fd_sc_hd__a21oi_2 _38559_ (.A1(_15683_),
    .A2(_15693_),
    .B1(_15686_),
    .Y(_15985_));
 sky130_fd_sc_hd__o21ai_2 _38560_ (.A1(_15749_),
    .A2(_15985_),
    .B1(_15694_),
    .Y(_15986_));
 sky130_fd_sc_hd__a21o_1 _38561_ (.A1(_15973_),
    .A2(_15979_),
    .B1(_15980_),
    .X(_15987_));
 sky130_fd_sc_hd__o21a_1 _38562_ (.A1(_15802_),
    .A2(_15803_),
    .B1(_15807_),
    .X(_15988_));
 sky130_fd_sc_hd__a21oi_4 _38563_ (.A1(_15804_),
    .A2(_15988_),
    .B1(_15808_),
    .Y(_15989_));
 sky130_fd_sc_hd__nand3_4 _38564_ (.A(_15973_),
    .B(_15980_),
    .C(_15979_),
    .Y(_15990_));
 sky130_fd_sc_hd__nand3_2 _38565_ (.A(_15987_),
    .B(_15989_),
    .C(_15990_),
    .Y(_15991_));
 sky130_fd_sc_hd__nand3_4 _38566_ (.A(_15984_),
    .B(_15986_),
    .C(_15991_),
    .Y(_15992_));
 sky130_fd_sc_hd__o21ai_2 _38567_ (.A1(_15981_),
    .A2(_15983_),
    .B1(_15989_),
    .Y(_15993_));
 sky130_fd_sc_hd__a21boi_2 _38568_ (.A1(_15738_),
    .A2(_15702_),
    .B1_N(_15694_),
    .Y(_15994_));
 sky130_fd_sc_hd__o211ai_2 _38569_ (.A1(_15808_),
    .A2(_15806_),
    .B1(_15990_),
    .C1(_15987_),
    .Y(_15995_));
 sky130_fd_sc_hd__nand3_4 _38570_ (.A(_15993_),
    .B(_15994_),
    .C(_15995_),
    .Y(_15996_));
 sky130_fd_sc_hd__nand2_1 _38571_ (.A(_15720_),
    .B(_15728_),
    .Y(_15997_));
 sky130_fd_sc_hd__nand2_2 _38572_ (.A(_15997_),
    .B(_15726_),
    .Y(_15998_));
 sky130_vsdinv _38573_ (.A(_15998_),
    .Y(_15999_));
 sky130_fd_sc_hd__nor2_1 _38574_ (.A(_14353_),
    .B(_15999_),
    .Y(_16000_));
 sky130_fd_sc_hd__clkbuf_2 _38575_ (.A(_16000_),
    .X(_16001_));
 sky130_fd_sc_hd__nor2_2 _38576_ (.A(_14930_),
    .B(_15998_),
    .Y(_16002_));
 sky130_fd_sc_hd__o2bb2ai_2 _38577_ (.A1_N(_15992_),
    .A2_N(_15996_),
    .B1(_16001_),
    .B2(_16002_),
    .Y(_16003_));
 sky130_fd_sc_hd__nand2_1 _38578_ (.A(_15751_),
    .B(_15762_),
    .Y(_16004_));
 sky130_fd_sc_hd__nand2_1 _38579_ (.A(_16004_),
    .B(_15740_),
    .Y(_16005_));
 sky130_fd_sc_hd__nor2_2 _38580_ (.A(_16002_),
    .B(_16000_),
    .Y(_16006_));
 sky130_fd_sc_hd__nand3_2 _38581_ (.A(_15996_),
    .B(_15992_),
    .C(_16006_),
    .Y(_16007_));
 sky130_fd_sc_hd__nand3_4 _38582_ (.A(_16003_),
    .B(_16005_),
    .C(_16007_),
    .Y(_16008_));
 sky130_fd_sc_hd__nor2_1 _38583_ (.A(_15754_),
    .B(_15998_),
    .Y(_16009_));
 sky130_fd_sc_hd__nor2_1 _38584_ (.A(_14931_),
    .B(_15999_),
    .Y(_16010_));
 sky130_fd_sc_hd__o2bb2ai_2 _38585_ (.A1_N(_15992_),
    .A2_N(_15996_),
    .B1(_16009_),
    .B2(_16010_),
    .Y(_16011_));
 sky130_fd_sc_hd__a21boi_2 _38586_ (.A1(_15751_),
    .A2(_15762_),
    .B1_N(_15740_),
    .Y(_16012_));
 sky130_fd_sc_hd__nand3b_4 _38587_ (.A_N(_16006_),
    .B(_15996_),
    .C(_15992_),
    .Y(_16013_));
 sky130_fd_sc_hd__nand3_4 _38588_ (.A(_16011_),
    .B(_16012_),
    .C(_16013_),
    .Y(_16014_));
 sky130_fd_sc_hd__nand3_4 _38589_ (.A(_16008_),
    .B(_16014_),
    .C(_15503_),
    .Y(_16015_));
 sky130_vsdinv _38590_ (.A(_16015_),
    .Y(_16016_));
 sky130_fd_sc_hd__o2bb2ai_2 _38591_ (.A1_N(_16008_),
    .A2_N(_16014_),
    .B1(net412),
    .B2(_15502_),
    .Y(_16017_));
 sky130_fd_sc_hd__a21oi_2 _38592_ (.A1(_15761_),
    .A2(_15763_),
    .B1(_15760_),
    .Y(_16018_));
 sky130_fd_sc_hd__o21ai_2 _38593_ (.A1(_15476_),
    .A2(_16018_),
    .B1(_15764_),
    .Y(_16019_));
 sky130_fd_sc_hd__nand2_2 _38594_ (.A(_16017_),
    .B(_16019_),
    .Y(_16020_));
 sky130_fd_sc_hd__a21o_1 _38595_ (.A1(_16017_),
    .A2(_16015_),
    .B1(_16019_),
    .X(_16021_));
 sky130_fd_sc_hd__o21ai_1 _38596_ (.A1(_16016_),
    .A2(_16020_),
    .B1(_16021_),
    .Y(_16022_));
 sky130_fd_sc_hd__o21ai_1 _38597_ (.A1(_15776_),
    .A2(_15783_),
    .B1(_15775_),
    .Y(_16023_));
 sky130_fd_sc_hd__xnor2_1 _38598_ (.A(_16022_),
    .B(_16023_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _38599_ (.A(_15843_),
    .B(_15850_),
    .Y(_16024_));
 sky130_fd_sc_hd__nand2_1 _38600_ (.A(_16024_),
    .B(_15848_),
    .Y(_16025_));
 sky130_fd_sc_hd__nor2_8 _38601_ (.A(_15787_),
    .B(_15832_),
    .Y(_16026_));
 sky130_vsdinv _38602_ (.A(_15789_),
    .Y(_16027_));
 sky130_fd_sc_hd__o31ai_2 _38603_ (.A1(_15787_),
    .A2(_15790_),
    .A3(_15788_),
    .B1(_16027_),
    .Y(_16028_));
 sky130_fd_sc_hd__or2_1 _38604_ (.A(_16026_),
    .B(_16028_),
    .X(_16029_));
 sky130_fd_sc_hd__nand2_1 _38605_ (.A(_16028_),
    .B(_16026_),
    .Y(_16030_));
 sky130_fd_sc_hd__nand2_1 _38606_ (.A(_16029_),
    .B(_16030_),
    .Y(_16031_));
 sky130_fd_sc_hd__nand2_1 _38607_ (.A(_16031_),
    .B(_13679_),
    .Y(_16032_));
 sky130_fd_sc_hd__nand3_1 _38608_ (.A(_16029_),
    .B(_14014_),
    .C(_16030_),
    .Y(_16033_));
 sky130_fd_sc_hd__nand2_1 _38609_ (.A(_16032_),
    .B(_16033_),
    .Y(_16034_));
 sky130_fd_sc_hd__or2_2 _38610_ (.A(_16025_),
    .B(_16034_),
    .X(_16035_));
 sky130_fd_sc_hd__nand2_2 _38611_ (.A(_16034_),
    .B(_16025_),
    .Y(_16036_));
 sky130_fd_sc_hd__nand2_2 _38612_ (.A(_15800_),
    .B(_15798_),
    .Y(_16037_));
 sky130_fd_sc_hd__a21o_1 _38613_ (.A1(_16035_),
    .A2(_16036_),
    .B1(_16037_),
    .X(_16038_));
 sky130_vsdinv _38614_ (.A(_16038_),
    .Y(_16039_));
 sky130_fd_sc_hd__nand3_4 _38615_ (.A(_16035_),
    .B(_16037_),
    .C(_16036_),
    .Y(_16040_));
 sky130_vsdinv _38616_ (.A(_16040_),
    .Y(_16041_));
 sky130_fd_sc_hd__a21oi_4 _38617_ (.A1(_15901_),
    .A2(_15900_),
    .B1(_15947_),
    .Y(_16042_));
 sky130_fd_sc_hd__nand2_2 _38618_ (.A(_19859_),
    .B(_12109_),
    .Y(_16043_));
 sky130_fd_sc_hd__nand2_1 _38619_ (.A(_10918_),
    .B(_20091_),
    .Y(_16044_));
 sky130_fd_sc_hd__nor2_2 _38620_ (.A(_16043_),
    .B(_16044_),
    .Y(_16045_));
 sky130_fd_sc_hd__nand2_1 _38621_ (.A(_19867_),
    .B(_20088_),
    .Y(_16046_));
 sky130_fd_sc_hd__and2_1 _38622_ (.A(_16043_),
    .B(_16044_),
    .X(_16047_));
 sky130_fd_sc_hd__or3_4 _38623_ (.A(_16045_),
    .B(_16046_),
    .C(_16047_),
    .X(_16048_));
 sky130_fd_sc_hd__o21ai_2 _38624_ (.A1(_16045_),
    .A2(_16047_),
    .B1(_16046_),
    .Y(_16049_));
 sky130_fd_sc_hd__nand2_1 _38625_ (.A(_16048_),
    .B(_16049_),
    .Y(_16050_));
 sky130_fd_sc_hd__nor2_1 _38626_ (.A(_15854_),
    .B(_15856_),
    .Y(_16051_));
 sky130_fd_sc_hd__nor2_2 _38627_ (.A(_16051_),
    .B(_15864_),
    .Y(_16052_));
 sky130_fd_sc_hd__nand2_2 _38628_ (.A(_16050_),
    .B(_16052_),
    .Y(_16053_));
 sky130_fd_sc_hd__nand3b_4 _38629_ (.A_N(_16052_),
    .B(_16048_),
    .C(_16049_),
    .Y(_16054_));
 sky130_fd_sc_hd__nand2_1 _38630_ (.A(_16053_),
    .B(_16054_),
    .Y(_16055_));
 sky130_fd_sc_hd__nand2_4 _38631_ (.A(_10768_),
    .B(_11165_),
    .Y(_16056_));
 sky130_fd_sc_hd__a22o_1 _38632_ (.A1(_10935_),
    .A2(_12298_),
    .B1(_10945_),
    .B2(_10768_),
    .X(_16057_));
 sky130_fd_sc_hd__o2111a_1 _38633_ (.A1(_15871_),
    .A2(_16056_),
    .B1(_19879_),
    .C1(_20075_),
    .D1(_16057_),
    .X(_16058_));
 sky130_fd_sc_hd__clkbuf_4 _38634_ (.A(_10772_),
    .X(_16059_));
 sky130_fd_sc_hd__o21ai_1 _38635_ (.A1(_15871_),
    .A2(_16056_),
    .B1(_16057_),
    .Y(_16060_));
 sky130_fd_sc_hd__o21a_1 _38636_ (.A1(_07141_),
    .A2(_16059_),
    .B1(_16060_),
    .X(_16061_));
 sky130_fd_sc_hd__nor2_2 _38637_ (.A(_16058_),
    .B(_16061_),
    .Y(_16062_));
 sky130_fd_sc_hd__nand2_1 _38638_ (.A(_16055_),
    .B(_16062_),
    .Y(_16063_));
 sky130_vsdinv _38639_ (.A(_16062_),
    .Y(_16064_));
 sky130_fd_sc_hd__nand3_2 _38640_ (.A(_16053_),
    .B(_16054_),
    .C(_16064_),
    .Y(_16065_));
 sky130_fd_sc_hd__nand3b_4 _38641_ (.A_N(_16042_),
    .B(_16063_),
    .C(_16065_),
    .Y(_16066_));
 sky130_fd_sc_hd__nand2_2 _38642_ (.A(_16053_),
    .B(_16062_),
    .Y(_16067_));
 sky130_vsdinv _38643_ (.A(_16054_),
    .Y(_16068_));
 sky130_fd_sc_hd__nand2_1 _38644_ (.A(_16055_),
    .B(_16064_),
    .Y(_16069_));
 sky130_fd_sc_hd__o211ai_4 _38645_ (.A1(_16067_),
    .A2(_16068_),
    .B1(_16042_),
    .C1(_16069_),
    .Y(_16070_));
 sky130_fd_sc_hd__nand2_4 _38646_ (.A(_15882_),
    .B(_15879_),
    .Y(_16071_));
 sky130_fd_sc_hd__a21oi_4 _38647_ (.A1(_16066_),
    .A2(_16070_),
    .B1(_16071_),
    .Y(_16072_));
 sky130_vsdinv _38648_ (.A(_16071_),
    .Y(_16073_));
 sky130_fd_sc_hd__nand2_4 _38649_ (.A(_16066_),
    .B(_16070_),
    .Y(_16074_));
 sky130_fd_sc_hd__nor2_8 _38650_ (.A(_16073_),
    .B(_16074_),
    .Y(_16075_));
 sky130_fd_sc_hd__nand2_1 _38651_ (.A(_15597_),
    .B(_11078_),
    .Y(_16076_));
 sky130_fd_sc_hd__nand2_1 _38652_ (.A(_15594_),
    .B(_20102_),
    .Y(_16077_));
 sky130_fd_sc_hd__nor2_1 _38653_ (.A(_16076_),
    .B(_16077_),
    .Y(_16078_));
 sky130_fd_sc_hd__and2_1 _38654_ (.A(_16076_),
    .B(_16077_),
    .X(_16079_));
 sky130_fd_sc_hd__or4_4 _38655_ (.A(_08615_),
    .B(_09880_),
    .C(_16078_),
    .D(_16079_),
    .X(_16080_));
 sky130_fd_sc_hd__a2bb2o_2 _38656_ (.A1_N(_16078_),
    .A2_N(_16079_),
    .B1(_19856_),
    .B2(_20099_),
    .X(_16081_));
 sky130_fd_sc_hd__a21o_1 _38657_ (.A1(_15928_),
    .A2(_15930_),
    .B1(_15927_),
    .X(_16082_));
 sky130_fd_sc_hd__a21o_2 _38658_ (.A1(_16080_),
    .A2(_16081_),
    .B1(_16082_),
    .X(_16083_));
 sky130_fd_sc_hd__nand3_4 _38659_ (.A(_16080_),
    .B(_16082_),
    .C(_16081_),
    .Y(_16084_));
 sky130_fd_sc_hd__nand2_1 _38660_ (.A(_16083_),
    .B(_16084_),
    .Y(_16085_));
 sky130_fd_sc_hd__nand2_4 _38661_ (.A(_15893_),
    .B(_15891_),
    .Y(_16086_));
 sky130_vsdinv _38662_ (.A(_16086_),
    .Y(_16087_));
 sky130_fd_sc_hd__nand2_2 _38663_ (.A(_16085_),
    .B(_16087_),
    .Y(_16088_));
 sky130_fd_sc_hd__nand3_4 _38664_ (.A(_16083_),
    .B(_16086_),
    .C(_16084_),
    .Y(_16089_));
 sky130_fd_sc_hd__nand2_8 _38665_ (.A(_16088_),
    .B(_16089_),
    .Y(_16090_));
 sky130_fd_sc_hd__nand2_2 _38666_ (.A(_19845_),
    .B(_20109_),
    .Y(_16091_));
 sky130_vsdinv _38667_ (.A(net463),
    .Y(_16092_));
 sky130_fd_sc_hd__clkbuf_2 _38668_ (.A(_16092_),
    .X(_16093_));
 sky130_vsdinv _38669_ (.A(_09997_),
    .Y(_16094_));
 sky130_vsdinv _38670_ (.A(_10412_),
    .Y(_16095_));
 sky130_fd_sc_hd__o22a_1 _38671_ (.A1(_16094_),
    .A2(_12073_),
    .B1(_16095_),
    .B2(_10824_),
    .X(_16096_));
 sky130_fd_sc_hd__a31o_1 _38672_ (.A1(_20112_),
    .A2(_20116_),
    .A3(_16093_),
    .B1(_16096_),
    .X(_16097_));
 sky130_fd_sc_hd__nor2_4 _38673_ (.A(_16091_),
    .B(_16097_),
    .Y(_16098_));
 sky130_fd_sc_hd__and2_2 _38674_ (.A(_16097_),
    .B(_16091_),
    .X(_16099_));
 sky130_fd_sc_hd__nor2_4 _38675_ (.A(_16098_),
    .B(_16099_),
    .Y(_16100_));
 sky130_fd_sc_hd__and4_1 _38676_ (.A(_11096_),
    .B(_18695_),
    .C(_15907_),
    .D(_20124_),
    .X(_16101_));
 sky130_fd_sc_hd__clkbuf_2 _38677_ (.A(_15915_),
    .X(_16102_));
 sky130_fd_sc_hd__buf_2 _38678_ (.A(_16102_),
    .X(_16103_));
 sky130_fd_sc_hd__o22a_1 _38679_ (.A1(_20127_),
    .A2(_11276_),
    .B1(_16103_),
    .B2(_11457_),
    .X(_16104_));
 sky130_fd_sc_hd__nor2_2 _38680_ (.A(_16101_),
    .B(_16104_),
    .Y(_16105_));
 sky130_fd_sc_hd__nand3_4 _38681_ (.A(_16105_),
    .B(_19834_),
    .C(_20120_),
    .Y(_16106_));
 sky130_fd_sc_hd__clkbuf_4 _38682_ (.A(_19833_),
    .X(_16107_));
 sky130_fd_sc_hd__nand2_1 _38683_ (.A(_16107_),
    .B(_20120_),
    .Y(_16108_));
 sky130_fd_sc_hd__o21ai_2 _38684_ (.A1(_16101_),
    .A2(_16104_),
    .B1(_16108_),
    .Y(_16109_));
 sky130_fd_sc_hd__a21o_1 _38685_ (.A1(_15917_),
    .A2(_15913_),
    .B1(_15906_),
    .X(_16110_));
 sky130_fd_sc_hd__a21o_2 _38686_ (.A1(_16106_),
    .A2(_16109_),
    .B1(_16110_),
    .X(_16111_));
 sky130_fd_sc_hd__nand3_4 _38687_ (.A(_16106_),
    .B(_16109_),
    .C(_16110_),
    .Y(_16112_));
 sky130_fd_sc_hd__nand3_4 _38688_ (.A(_16100_),
    .B(_16111_),
    .C(_16112_),
    .Y(_16113_));
 sky130_fd_sc_hd__o2bb2ai_4 _38689_ (.A1_N(_16112_),
    .A2_N(_16111_),
    .B1(_16098_),
    .B2(_16099_),
    .Y(_16114_));
 sky130_fd_sc_hd__nand2_4 _38690_ (.A(_15943_),
    .B(_15919_),
    .Y(_16115_));
 sky130_fd_sc_hd__nand3_4 _38691_ (.A(_16113_),
    .B(_16114_),
    .C(_16115_),
    .Y(_16116_));
 sky130_fd_sc_hd__a21o_1 _38692_ (.A1(_16113_),
    .A2(_16114_),
    .B1(_16115_),
    .X(_16117_));
 sky130_fd_sc_hd__nand3b_4 _38693_ (.A_N(_16090_),
    .B(_16116_),
    .C(_16117_),
    .Y(_16118_));
 sky130_fd_sc_hd__a21oi_4 _38694_ (.A1(_16113_),
    .A2(_16114_),
    .B1(_16115_),
    .Y(_16119_));
 sky130_fd_sc_hd__and3_1 _38695_ (.A(_16113_),
    .B(_16114_),
    .C(_16115_),
    .X(_16120_));
 sky130_fd_sc_hd__o21ai_4 _38696_ (.A1(_16119_),
    .A2(_16120_),
    .B1(_16090_),
    .Y(_16121_));
 sky130_fd_sc_hd__and2_2 _38697_ (.A(_15946_),
    .B(_15951_),
    .X(_16122_));
 sky130_fd_sc_hd__nor2_4 _38698_ (.A(_15944_),
    .B(_16122_),
    .Y(_16123_));
 sky130_fd_sc_hd__a21boi_4 _38699_ (.A1(_16118_),
    .A2(_16121_),
    .B1_N(_16123_),
    .Y(_16124_));
 sky130_fd_sc_hd__o211a_1 _38700_ (.A1(_15944_),
    .A2(_16122_),
    .B1(_16121_),
    .C1(_16118_),
    .X(_16125_));
 sky130_fd_sc_hd__o22ai_4 _38701_ (.A1(_16072_),
    .A2(_16075_),
    .B1(_16124_),
    .B2(_16125_),
    .Y(_16126_));
 sky130_fd_sc_hd__nand2_1 _38702_ (.A(_15961_),
    .B(_15962_),
    .Y(_16127_));
 sky130_fd_sc_hd__nand2_4 _38703_ (.A(_16127_),
    .B(_15963_),
    .Y(_16128_));
 sky130_fd_sc_hd__nand2_1 _38704_ (.A(_16118_),
    .B(_16121_),
    .Y(_16129_));
 sky130_fd_sc_hd__nand2_4 _38705_ (.A(_16129_),
    .B(_16123_),
    .Y(_16130_));
 sky130_fd_sc_hd__nand2_1 _38706_ (.A(_16117_),
    .B(_16116_),
    .Y(_16131_));
 sky130_fd_sc_hd__a21oi_4 _38707_ (.A1(_16131_),
    .A2(_16090_),
    .B1(_16123_),
    .Y(_16132_));
 sky130_fd_sc_hd__nand2_4 _38708_ (.A(_16132_),
    .B(_16118_),
    .Y(_16133_));
 sky130_fd_sc_hd__nor2_8 _38709_ (.A(_16072_),
    .B(_16075_),
    .Y(_16134_));
 sky130_fd_sc_hd__nand3_4 _38710_ (.A(_16130_),
    .B(_16133_),
    .C(_16134_),
    .Y(_16135_));
 sky130_fd_sc_hd__nand3_4 _38711_ (.A(_16126_),
    .B(_16128_),
    .C(_16135_),
    .Y(_16136_));
 sky130_fd_sc_hd__o21ai_2 _38712_ (.A1(_16124_),
    .A2(_16125_),
    .B1(_16134_),
    .Y(_16137_));
 sky130_fd_sc_hd__a21o_1 _38713_ (.A1(_15879_),
    .A2(_15882_),
    .B1(_16074_),
    .X(_16138_));
 sky130_fd_sc_hd__nand2_1 _38714_ (.A(_16074_),
    .B(_16073_),
    .Y(_16139_));
 sky130_fd_sc_hd__nand2_2 _38715_ (.A(_16138_),
    .B(_16139_),
    .Y(_16140_));
 sky130_fd_sc_hd__nand3_4 _38716_ (.A(_16130_),
    .B(_16133_),
    .C(_16140_),
    .Y(_16141_));
 sky130_vsdinv _38717_ (.A(_16128_),
    .Y(_16142_));
 sky130_fd_sc_hd__nand3_4 _38718_ (.A(_16137_),
    .B(_16141_),
    .C(_16142_),
    .Y(_16143_));
 sky130_fd_sc_hd__a21boi_4 _38719_ (.A1(_15881_),
    .A2(_15886_),
    .B1_N(_15884_),
    .Y(_16144_));
 sky130_fd_sc_hd__o21ba_4 _38720_ (.A1(_15871_),
    .A2(_15867_),
    .B1_N(_15870_),
    .X(_16145_));
 sky130_vsdinv _38721_ (.A(_07294_),
    .Y(_16146_));
 sky130_fd_sc_hd__clkbuf_4 _38722_ (.A(_11176_),
    .X(_16147_));
 sky130_fd_sc_hd__nand2_4 _38723_ (.A(_11975_),
    .B(_07291_),
    .Y(_16148_));
 sky130_fd_sc_hd__o21ai_4 _38724_ (.A1(_16146_),
    .A2(_16147_),
    .B1(_16148_),
    .Y(_16149_));
 sky130_fd_sc_hd__or3_4 _38725_ (.A(_16148_),
    .B(_16146_),
    .C(_11176_),
    .X(_16150_));
 sky130_fd_sc_hd__o2bb2ai_4 _38726_ (.A1_N(_16149_),
    .A2_N(_16150_),
    .B1(_13024_),
    .B2(net443),
    .Y(_16151_));
 sky130_fd_sc_hd__nand3_4 _38727_ (.A(_16150_),
    .B(_15816_),
    .C(_16149_),
    .Y(_16152_));
 sky130_fd_sc_hd__nand2_4 _38728_ (.A(_16151_),
    .B(_16152_),
    .Y(_16153_));
 sky130_fd_sc_hd__nor2_8 _38729_ (.A(_16145_),
    .B(_16153_),
    .Y(_16154_));
 sky130_fd_sc_hd__nand2_4 _38730_ (.A(_15818_),
    .B(_15815_),
    .Y(_16155_));
 sky130_fd_sc_hd__nand2_4 _38731_ (.A(_16153_),
    .B(_16145_),
    .Y(_16156_));
 sky130_fd_sc_hd__nand3b_2 _38732_ (.A_N(_16154_),
    .B(_16155_),
    .C(_16156_),
    .Y(_16157_));
 sky130_fd_sc_hd__nand2_2 _38733_ (.A(_15824_),
    .B(_15821_),
    .Y(_16158_));
 sky130_vsdinv _38734_ (.A(_15871_),
    .Y(_16159_));
 sky130_fd_sc_hd__a31o_1 _38735_ (.A1(_20084_),
    .A2(_20089_),
    .A3(_16159_),
    .B1(_15870_),
    .X(_16160_));
 sky130_fd_sc_hd__a21oi_4 _38736_ (.A1(_16151_),
    .A2(_16152_),
    .B1(_16160_),
    .Y(_16161_));
 sky130_vsdinv _38737_ (.A(_16155_),
    .Y(_16162_));
 sky130_fd_sc_hd__o21ai_2 _38738_ (.A1(_16161_),
    .A2(_16154_),
    .B1(_16162_),
    .Y(_16163_));
 sky130_fd_sc_hd__nand3_4 _38739_ (.A(_16157_),
    .B(_16158_),
    .C(_16163_),
    .Y(_16164_));
 sky130_fd_sc_hd__nand3b_2 _38740_ (.A_N(_16154_),
    .B(_16162_),
    .C(_16156_),
    .Y(_16165_));
 sky130_vsdinv _38741_ (.A(_16158_),
    .Y(_16166_));
 sky130_fd_sc_hd__o21ai_2 _38742_ (.A1(_16161_),
    .A2(_16154_),
    .B1(_16155_),
    .Y(_16167_));
 sky130_fd_sc_hd__nand3_4 _38743_ (.A(_16165_),
    .B(_16166_),
    .C(_16167_),
    .Y(_16168_));
 sky130_fd_sc_hd__nand2_1 _38744_ (.A(_16164_),
    .B(_16168_),
    .Y(_16169_));
 sky130_fd_sc_hd__clkbuf_4 _38745_ (.A(_15840_),
    .X(_16170_));
 sky130_fd_sc_hd__nand2_1 _38746_ (.A(_16169_),
    .B(_16170_),
    .Y(_16171_));
 sky130_fd_sc_hd__clkbuf_4 _38747_ (.A(_15835_),
    .X(_16172_));
 sky130_fd_sc_hd__nand3_2 _38748_ (.A(_16164_),
    .B(_16168_),
    .C(_16172_),
    .Y(_16173_));
 sky130_fd_sc_hd__nand3b_4 _38749_ (.A_N(_16144_),
    .B(_16171_),
    .C(_16173_),
    .Y(_16174_));
 sky130_fd_sc_hd__nand2_1 _38750_ (.A(_16169_),
    .B(_16172_),
    .Y(_16175_));
 sky130_fd_sc_hd__nand3_2 _38751_ (.A(_16164_),
    .B(_16168_),
    .C(_16170_),
    .Y(_16176_));
 sky130_fd_sc_hd__nand3_4 _38752_ (.A(_16175_),
    .B(_16144_),
    .C(_16176_),
    .Y(_16177_));
 sky130_fd_sc_hd__nor2_2 _38753_ (.A(_15830_),
    .B(_16170_),
    .Y(_16178_));
 sky130_fd_sc_hd__nor2_4 _38754_ (.A(_15827_),
    .B(_16178_),
    .Y(_16179_));
 sky130_vsdinv _38755_ (.A(_16179_),
    .Y(_16180_));
 sky130_fd_sc_hd__a21oi_4 _38756_ (.A1(_16174_),
    .A2(_16177_),
    .B1(_16180_),
    .Y(_16181_));
 sky130_fd_sc_hd__nand2_2 _38757_ (.A(_16174_),
    .B(_16177_),
    .Y(_16182_));
 sky130_fd_sc_hd__nor2_4 _38758_ (.A(_16179_),
    .B(_16182_),
    .Y(_16183_));
 sky130_fd_sc_hd__o2bb2ai_4 _38759_ (.A1_N(_16136_),
    .A2_N(_16143_),
    .B1(_16181_),
    .B2(_16183_),
    .Y(_16184_));
 sky130_fd_sc_hd__nor2_4 _38760_ (.A(_16181_),
    .B(_16183_),
    .Y(_16185_));
 sky130_fd_sc_hd__nand3_4 _38761_ (.A(_16185_),
    .B(_16143_),
    .C(_16136_),
    .Y(_16186_));
 sky130_fd_sc_hd__nand2_4 _38762_ (.A(_15979_),
    .B(_15978_),
    .Y(_16187_));
 sky130_fd_sc_hd__a21oi_4 _38763_ (.A1(_16184_),
    .A2(_16186_),
    .B1(_16187_),
    .Y(_16188_));
 sky130_fd_sc_hd__and3_1 _38764_ (.A(_16126_),
    .B(_16128_),
    .C(_16135_),
    .X(_16189_));
 sky130_fd_sc_hd__nand2_2 _38765_ (.A(_16185_),
    .B(_16143_),
    .Y(_16190_));
 sky130_fd_sc_hd__o211a_1 _38766_ (.A1(_16189_),
    .A2(_16190_),
    .B1(_16187_),
    .C1(_16184_),
    .X(_16191_));
 sky130_fd_sc_hd__o22ai_4 _38767_ (.A1(_16039_),
    .A2(_16041_),
    .B1(_16188_),
    .B2(_16191_),
    .Y(_16192_));
 sky130_fd_sc_hd__nand2_2 _38768_ (.A(_16038_),
    .B(_16040_),
    .Y(_16193_));
 sky130_fd_sc_hd__nand2_1 _38769_ (.A(_16184_),
    .B(_16186_),
    .Y(_16194_));
 sky130_vsdinv _38770_ (.A(_16187_),
    .Y(_16195_));
 sky130_fd_sc_hd__nand2_2 _38771_ (.A(_16194_),
    .B(_16195_),
    .Y(_16196_));
 sky130_fd_sc_hd__nand3_4 _38772_ (.A(_16184_),
    .B(_16187_),
    .C(_16186_),
    .Y(_16197_));
 sky130_fd_sc_hd__nand3b_4 _38773_ (.A_N(_16193_),
    .B(_16196_),
    .C(_16197_),
    .Y(_16198_));
 sky130_fd_sc_hd__nand2_1 _38774_ (.A(_15987_),
    .B(_15989_),
    .Y(_16199_));
 sky130_fd_sc_hd__nand2_4 _38775_ (.A(_16199_),
    .B(_15990_),
    .Y(_16200_));
 sky130_fd_sc_hd__a21oi_4 _38776_ (.A1(_16192_),
    .A2(_16198_),
    .B1(_16200_),
    .Y(_16201_));
 sky130_fd_sc_hd__and3_2 _38777_ (.A(_16192_),
    .B(_16198_),
    .C(_16200_),
    .X(_16202_));
 sky130_fd_sc_hd__nand2_1 _38778_ (.A(_15988_),
    .B(_15804_),
    .Y(_16203_));
 sky130_fd_sc_hd__and2_2 _38779_ (.A(_16203_),
    .B(_15801_),
    .X(_16204_));
 sky130_fd_sc_hd__nor2_8 _38780_ (.A(_14353_),
    .B(_16204_),
    .Y(_16205_));
 sky130_vsdinv _38781_ (.A(_16205_),
    .Y(_16206_));
 sky130_fd_sc_hd__nand2_1 _38782_ (.A(_16204_),
    .B(_14354_),
    .Y(_16207_));
 sky130_fd_sc_hd__nand2_2 _38783_ (.A(_16206_),
    .B(_16207_),
    .Y(_16208_));
 sky130_fd_sc_hd__o21ai_1 _38784_ (.A1(_16201_),
    .A2(_16202_),
    .B1(_16208_),
    .Y(_16209_));
 sky130_fd_sc_hd__nand2_1 _38785_ (.A(_15996_),
    .B(_16006_),
    .Y(_16210_));
 sky130_fd_sc_hd__nand2_1 _38786_ (.A(_16210_),
    .B(_15992_),
    .Y(_16211_));
 sky130_fd_sc_hd__a21o_2 _38787_ (.A1(_16192_),
    .A2(_16198_),
    .B1(_16200_),
    .X(_16212_));
 sky130_fd_sc_hd__nand3_4 _38788_ (.A(_16192_),
    .B(_16198_),
    .C(_16200_),
    .Y(_16213_));
 sky130_vsdinv _38789_ (.A(_16208_),
    .Y(_16214_));
 sky130_fd_sc_hd__nand3_1 _38790_ (.A(_16212_),
    .B(_16213_),
    .C(_16214_),
    .Y(_16215_));
 sky130_fd_sc_hd__nand3_2 _38791_ (.A(_16209_),
    .B(_16211_),
    .C(_16215_),
    .Y(_16216_));
 sky130_fd_sc_hd__o21ai_4 _38792_ (.A1(_16201_),
    .A2(_16202_),
    .B1(_16214_),
    .Y(_16217_));
 sky130_vsdinv _38793_ (.A(_16211_),
    .Y(_16218_));
 sky130_fd_sc_hd__nand3_4 _38794_ (.A(_16212_),
    .B(_16213_),
    .C(_16208_),
    .Y(_16219_));
 sky130_fd_sc_hd__nand3_4 _38795_ (.A(_16217_),
    .B(_16218_),
    .C(_16219_),
    .Y(_16220_));
 sky130_fd_sc_hd__a21oi_2 _38796_ (.A1(_16216_),
    .A2(_16220_),
    .B1(_16001_),
    .Y(_16221_));
 sky130_fd_sc_hd__and3_1 _38797_ (.A(_16216_),
    .B(_16220_),
    .C(_16001_),
    .X(_16222_));
 sky130_fd_sc_hd__a21bo_1 _38798_ (.A1(_15503_),
    .A2(_16014_),
    .B1_N(_16008_),
    .X(_16223_));
 sky130_fd_sc_hd__o21bai_4 _38799_ (.A1(_16221_),
    .A2(_16222_),
    .B1_N(_16223_),
    .Y(_16224_));
 sky130_fd_sc_hd__a21oi_4 _38800_ (.A1(_16217_),
    .A2(_16219_),
    .B1(_16218_),
    .Y(_16225_));
 sky130_fd_sc_hd__nand2_1 _38801_ (.A(_16220_),
    .B(_16001_),
    .Y(_16226_));
 sky130_fd_sc_hd__a21o_1 _38802_ (.A1(_16216_),
    .A2(_16220_),
    .B1(_16001_),
    .X(_16227_));
 sky130_fd_sc_hd__o211ai_4 _38803_ (.A1(_16225_),
    .A2(_16226_),
    .B1(_16223_),
    .C1(_16227_),
    .Y(_16228_));
 sky130_fd_sc_hd__nand2_1 _38804_ (.A(_16224_),
    .B(_16228_),
    .Y(_16229_));
 sky130_fd_sc_hd__nor3_4 _38805_ (.A(_14667_),
    .B(_15226_),
    .C(_14049_),
    .Y(_16230_));
 sky130_fd_sc_hd__o2111ai_4 _38806_ (.A1(_16016_),
    .A2(_16020_),
    .B1(_15775_),
    .C1(_15772_),
    .D1(_16021_),
    .Y(_16231_));
 sky130_fd_sc_hd__nor2_1 _38807_ (.A(_16231_),
    .B(_15780_),
    .Y(_16232_));
 sky130_fd_sc_hd__nand2_1 _38808_ (.A(_16230_),
    .B(_16232_),
    .Y(_16233_));
 sky130_fd_sc_hd__a21oi_1 _38809_ (.A1(_16017_),
    .A2(_16015_),
    .B1(_16019_),
    .Y(_16234_));
 sky130_fd_sc_hd__o22a_1 _38810_ (.A1(_16016_),
    .A2(_16020_),
    .B1(_15775_),
    .B2(_16234_),
    .X(_16235_));
 sky130_fd_sc_hd__o21ai_1 _38811_ (.A1(_16231_),
    .A2(_15782_),
    .B1(_16235_),
    .Y(_16236_));
 sky130_fd_sc_hd__a21oi_1 _38812_ (.A1(_15232_),
    .A2(_16232_),
    .B1(_16236_),
    .Y(_16237_));
 sky130_fd_sc_hd__o21a_4 _38813_ (.A1(_14055_),
    .A2(_16233_),
    .B1(_16237_),
    .X(_16238_));
 sky130_fd_sc_hd__nand3b_2 _38814_ (.A_N(_16231_),
    .B(_15225_),
    .C(_15497_),
    .Y(_16239_));
 sky130_fd_sc_hd__nor2_2 _38815_ (.A(_16239_),
    .B(_15228_),
    .Y(_16240_));
 sky130_fd_sc_hd__nand3_4 _38816_ (.A(net409),
    .B(_14052_),
    .C(_16240_),
    .Y(_16241_));
 sky130_fd_sc_hd__nand2_2 _38817_ (.A(_16238_),
    .B(_16241_),
    .Y(_16242_));
 sky130_fd_sc_hd__xnor2_1 _38818_ (.A(_16229_),
    .B(_16242_),
    .Y(_02667_));
 sky130_vsdinv _38819_ (.A(_16001_),
    .Y(_16243_));
 sky130_fd_sc_hd__a31oi_4 _38820_ (.A1(_16217_),
    .A2(_16218_),
    .A3(_16219_),
    .B1(_16243_),
    .Y(_16244_));
 sky130_fd_sc_hd__nor2_2 _38821_ (.A(_16225_),
    .B(_16244_),
    .Y(_16245_));
 sky130_fd_sc_hd__a21oi_4 _38822_ (.A1(_16212_),
    .A2(_16214_),
    .B1(_16202_),
    .Y(_16246_));
 sky130_fd_sc_hd__nand2_4 _38823_ (.A(_16040_),
    .B(_16036_),
    .Y(_16247_));
 sky130_fd_sc_hd__and2_2 _38824_ (.A(_16247_),
    .B(_15754_),
    .X(_16248_));
 sky130_fd_sc_hd__nor2_4 _38825_ (.A(_14354_),
    .B(_16247_),
    .Y(_16249_));
 sky130_fd_sc_hd__nand2_1 _38826_ (.A(_16197_),
    .B(_16193_),
    .Y(_16250_));
 sky130_fd_sc_hd__nand2_2 _38827_ (.A(_16177_),
    .B(_16180_),
    .Y(_16251_));
 sky130_fd_sc_hd__nor2_8 _38828_ (.A(_16027_),
    .B(_16026_),
    .Y(_16252_));
 sky130_fd_sc_hd__and2_2 _38829_ (.A(_16026_),
    .B(_15790_),
    .X(_16253_));
 sky130_fd_sc_hd__o21a_1 _38830_ (.A1(_16252_),
    .A2(_16253_),
    .B1(_13678_),
    .X(_16254_));
 sky130_fd_sc_hd__nor3_4 _38831_ (.A(_16253_),
    .B(_16252_),
    .C(_13678_),
    .Y(_16255_));
 sky130_fd_sc_hd__nor2_4 _38832_ (.A(_16254_),
    .B(_16255_),
    .Y(_16256_));
 sky130_vsdinv _38833_ (.A(_16256_),
    .Y(_16257_));
 sky130_fd_sc_hd__clkbuf_4 _38834_ (.A(_16257_),
    .X(_16258_));
 sky130_fd_sc_hd__a21o_1 _38835_ (.A1(_16251_),
    .A2(_16174_),
    .B1(_16258_),
    .X(_16259_));
 sky130_fd_sc_hd__nand3_2 _38836_ (.A(_16251_),
    .B(_16258_),
    .C(_16174_),
    .Y(_16260_));
 sky130_fd_sc_hd__nand2_1 _38837_ (.A(_16259_),
    .B(_16260_),
    .Y(_16261_));
 sky130_fd_sc_hd__and2_1 _38838_ (.A(_16031_),
    .B(_14014_),
    .X(_16262_));
 sky130_fd_sc_hd__nor2_1 _38839_ (.A(_16252_),
    .B(_16262_),
    .Y(_16263_));
 sky130_fd_sc_hd__nand2_1 _38840_ (.A(_16261_),
    .B(_16263_),
    .Y(_16264_));
 sky130_vsdinv _38841_ (.A(_16264_),
    .Y(_16265_));
 sky130_vsdinv _38842_ (.A(_16263_),
    .Y(_16266_));
 sky130_fd_sc_hd__and3_2 _38843_ (.A(_16266_),
    .B(_16259_),
    .C(_16260_),
    .X(_16267_));
 sky130_vsdinv _38844_ (.A(_16045_),
    .Y(_16268_));
 sky130_fd_sc_hd__and2_1 _38845_ (.A(_16048_),
    .B(_16268_),
    .X(_16269_));
 sky130_fd_sc_hd__nand2_1 _38846_ (.A(_11396_),
    .B(_11927_),
    .Y(_16270_));
 sky130_fd_sc_hd__nand2_1 _38847_ (.A(_12855_),
    .B(_10262_),
    .Y(_16271_));
 sky130_fd_sc_hd__or2_2 _38848_ (.A(_16270_),
    .B(_16271_),
    .X(_16272_));
 sky130_fd_sc_hd__nand2_1 _38849_ (.A(_16270_),
    .B(_16271_),
    .Y(_16273_));
 sky130_fd_sc_hd__nor2_2 _38850_ (.A(_07822_),
    .B(_10763_),
    .Y(_16274_));
 sky130_fd_sc_hd__a21o_1 _38851_ (.A1(_16272_),
    .A2(_16273_),
    .B1(_16274_),
    .X(_16275_));
 sky130_fd_sc_hd__nand3_2 _38852_ (.A(_16272_),
    .B(_16273_),
    .C(_16274_),
    .Y(_16276_));
 sky130_fd_sc_hd__nand2_1 _38853_ (.A(_16275_),
    .B(_16276_),
    .Y(_16277_));
 sky130_fd_sc_hd__nand2_2 _38854_ (.A(_16269_),
    .B(_16277_),
    .Y(_16278_));
 sky130_fd_sc_hd__a21o_1 _38855_ (.A1(_16268_),
    .A2(_16048_),
    .B1(_16277_),
    .X(_16279_));
 sky130_fd_sc_hd__nand2_1 _38856_ (.A(_19879_),
    .B(_10779_),
    .Y(_16280_));
 sky130_fd_sc_hd__nand2_2 _38857_ (.A(_11607_),
    .B(_13647_),
    .Y(_16281_));
 sky130_fd_sc_hd__a22o_1 _38858_ (.A1(_19871_),
    .A2(_20079_),
    .B1(_19875_),
    .B2(_20074_),
    .X(_16282_));
 sky130_fd_sc_hd__o21ai_1 _38859_ (.A1(_15871_),
    .A2(_16281_),
    .B1(_16282_),
    .Y(_16283_));
 sky130_fd_sc_hd__nor2_1 _38860_ (.A(_16280_),
    .B(_16283_),
    .Y(_16284_));
 sky130_fd_sc_hd__and2_1 _38861_ (.A(_16283_),
    .B(_16280_),
    .X(_16285_));
 sky130_fd_sc_hd__or2_4 _38862_ (.A(_16284_),
    .B(_16285_),
    .X(_16286_));
 sky130_fd_sc_hd__a21oi_2 _38863_ (.A1(_16278_),
    .A2(_16279_),
    .B1(_16286_),
    .Y(_16287_));
 sky130_fd_sc_hd__nand3_4 _38864_ (.A(_16278_),
    .B(_16279_),
    .C(_16286_),
    .Y(_16288_));
 sky130_vsdinv _38865_ (.A(_16288_),
    .Y(_16289_));
 sky130_fd_sc_hd__a21boi_4 _38866_ (.A1(_16083_),
    .A2(_16086_),
    .B1_N(_16084_),
    .Y(_16290_));
 sky130_fd_sc_hd__o21bai_4 _38867_ (.A1(_16287_),
    .A2(_16289_),
    .B1_N(_16290_),
    .Y(_16291_));
 sky130_fd_sc_hd__a21o_2 _38868_ (.A1(_16278_),
    .A2(_16279_),
    .B1(_16286_),
    .X(_16292_));
 sky130_fd_sc_hd__nand3_4 _38869_ (.A(_16292_),
    .B(_16290_),
    .C(_16288_),
    .Y(_16293_));
 sky130_fd_sc_hd__nand2_2 _38870_ (.A(_16067_),
    .B(_16054_),
    .Y(_16294_));
 sky130_fd_sc_hd__a21oi_4 _38871_ (.A1(_16291_),
    .A2(_16293_),
    .B1(_16294_),
    .Y(_16295_));
 sky130_vsdinv _38872_ (.A(_16294_),
    .Y(_16296_));
 sky130_fd_sc_hd__a31oi_4 _38873_ (.A1(_16292_),
    .A2(_16290_),
    .A3(_16288_),
    .B1(_16296_),
    .Y(_16297_));
 sky130_fd_sc_hd__nand2_1 _38874_ (.A(_16297_),
    .B(_16291_),
    .Y(_16298_));
 sky130_vsdinv _38875_ (.A(_16298_),
    .Y(_16299_));
 sky130_fd_sc_hd__a21boi_4 _38876_ (.A1(_16100_),
    .A2(_16111_),
    .B1_N(_16112_),
    .Y(_16300_));
 sky130_fd_sc_hd__and4_1 _38877_ (.A(_11457_),
    .B(_18695_),
    .C(_15907_),
    .D(_20120_),
    .X(_16301_));
 sky130_fd_sc_hd__o22a_2 _38878_ (.A1(_20124_),
    .A2(_15914_),
    .B1(_16103_),
    .B2(_10704_),
    .X(_16302_));
 sky130_fd_sc_hd__a211o_2 _38879_ (.A1(_19834_),
    .A2(_20116_),
    .B1(_16301_),
    .C1(_16302_),
    .X(_16303_));
 sky130_fd_sc_hd__nand2_1 _38880_ (.A(_16107_),
    .B(_20116_),
    .Y(_16304_));
 sky130_fd_sc_hd__o21bai_4 _38881_ (.A1(_16301_),
    .A2(_16302_),
    .B1_N(_16304_),
    .Y(_16305_));
 sky130_fd_sc_hd__o21ba_2 _38882_ (.A1(_16108_),
    .A2(_16104_),
    .B1_N(_16101_),
    .X(_16306_));
 sky130_fd_sc_hd__a21o_1 _38883_ (.A1(_16303_),
    .A2(_16305_),
    .B1(_16306_),
    .X(_16307_));
 sky130_fd_sc_hd__nand3_4 _38884_ (.A(_16303_),
    .B(_16305_),
    .C(_16306_),
    .Y(_16308_));
 sky130_fd_sc_hd__nand2_1 _38885_ (.A(_19844_),
    .B(_20106_),
    .Y(_16309_));
 sky130_vsdinv _38886_ (.A(_16309_),
    .Y(_16310_));
 sky130_fd_sc_hd__buf_4 _38887_ (.A(net440),
    .X(_16311_));
 sky130_fd_sc_hd__a22o_1 _38888_ (.A1(_15924_),
    .A2(_20112_),
    .B1(_19842_),
    .B2(_20109_),
    .X(_16312_));
 sky130_fd_sc_hd__o31ai_4 _38889_ (.A1(_16311_),
    .A2(_12093_),
    .A3(_15929_),
    .B1(_16312_),
    .Y(_16313_));
 sky130_fd_sc_hd__xor2_4 _38890_ (.A(_16310_),
    .B(_16313_),
    .X(_16314_));
 sky130_fd_sc_hd__a21o_4 _38891_ (.A1(_16307_),
    .A2(_16308_),
    .B1(_16314_),
    .X(_16315_));
 sky130_fd_sc_hd__nand3_4 _38892_ (.A(_16307_),
    .B(_16308_),
    .C(_16314_),
    .Y(_16316_));
 sky130_fd_sc_hd__nand3_4 _38893_ (.A(_16300_),
    .B(_16315_),
    .C(_16316_),
    .Y(_16317_));
 sky130_fd_sc_hd__a21o_1 _38894_ (.A1(_16315_),
    .A2(_16316_),
    .B1(_16300_),
    .X(_16318_));
 sky130_fd_sc_hd__nor2_1 _38895_ (.A(_08615_),
    .B(_11563_),
    .Y(_16319_));
 sky130_fd_sc_hd__nand2_1 _38896_ (.A(_15597_),
    .B(_20102_),
    .Y(_16320_));
 sky130_fd_sc_hd__nand2_1 _38897_ (.A(_15594_),
    .B(_20098_),
    .Y(_16321_));
 sky130_fd_sc_hd__nor2_2 _38898_ (.A(_16320_),
    .B(_16321_),
    .Y(_16322_));
 sky130_fd_sc_hd__and2_1 _38899_ (.A(_16320_),
    .B(_16321_),
    .X(_16323_));
 sky130_fd_sc_hd__nor2_1 _38900_ (.A(_16322_),
    .B(_16323_),
    .Y(_16324_));
 sky130_fd_sc_hd__or2_2 _38901_ (.A(_16319_),
    .B(_16324_),
    .X(_16325_));
 sky130_fd_sc_hd__nand2_2 _38902_ (.A(_16324_),
    .B(_16319_),
    .Y(_16326_));
 sky130_fd_sc_hd__buf_6 _38903_ (.A(_16311_),
    .X(_16327_));
 sky130_fd_sc_hd__o32ai_4 _38904_ (.A1(_15929_),
    .A2(_11074_),
    .A3(_16327_),
    .B1(_16091_),
    .B2(_16096_),
    .Y(_16328_));
 sky130_fd_sc_hd__a21o_1 _38905_ (.A1(_16325_),
    .A2(_16326_),
    .B1(_16328_),
    .X(_16329_));
 sky130_fd_sc_hd__o21ai_2 _38906_ (.A1(_16076_),
    .A2(_16077_),
    .B1(_16080_),
    .Y(_16330_));
 sky130_fd_sc_hd__nand3_4 _38907_ (.A(_16325_),
    .B(_16328_),
    .C(_16326_),
    .Y(_16331_));
 sky130_fd_sc_hd__nand3_2 _38908_ (.A(_16329_),
    .B(_16330_),
    .C(_16331_),
    .Y(_16332_));
 sky130_vsdinv _38909_ (.A(_16332_),
    .Y(_16333_));
 sky130_fd_sc_hd__nand2_1 _38910_ (.A(_16329_),
    .B(_16331_),
    .Y(_16334_));
 sky130_vsdinv _38911_ (.A(_16330_),
    .Y(_16335_));
 sky130_fd_sc_hd__nand2_1 _38912_ (.A(_16334_),
    .B(_16335_),
    .Y(_16336_));
 sky130_vsdinv _38913_ (.A(_16336_),
    .Y(_16337_));
 sky130_fd_sc_hd__o2bb2ai_4 _38914_ (.A1_N(_16317_),
    .A2_N(_16318_),
    .B1(_16333_),
    .B2(_16337_),
    .Y(_16338_));
 sky130_fd_sc_hd__and2_2 _38915_ (.A(_16336_),
    .B(_16332_),
    .X(_16339_));
 sky130_fd_sc_hd__nand3_4 _38916_ (.A(_16339_),
    .B(_16318_),
    .C(_16317_),
    .Y(_16340_));
 sky130_fd_sc_hd__o21ai_4 _38917_ (.A1(_16119_),
    .A2(_16090_),
    .B1(_16116_),
    .Y(_16341_));
 sky130_fd_sc_hd__a21oi_4 _38918_ (.A1(_16338_),
    .A2(_16340_),
    .B1(_16341_),
    .Y(_16342_));
 sky130_fd_sc_hd__nor2_1 _38919_ (.A(_16119_),
    .B(_16090_),
    .Y(_16343_));
 sky130_fd_sc_hd__o211a_4 _38920_ (.A1(_16120_),
    .A2(_16343_),
    .B1(_16340_),
    .C1(_16338_),
    .X(_16344_));
 sky130_fd_sc_hd__o22ai_4 _38921_ (.A1(_16295_),
    .A2(_16299_),
    .B1(_16342_),
    .B2(_16344_),
    .Y(_16345_));
 sky130_fd_sc_hd__o21ai_2 _38922_ (.A1(_16140_),
    .A2(_16124_),
    .B1(_16133_),
    .Y(_16346_));
 sky130_fd_sc_hd__a21o_2 _38923_ (.A1(_16338_),
    .A2(_16340_),
    .B1(_16341_),
    .X(_16347_));
 sky130_fd_sc_hd__a21oi_4 _38924_ (.A1(_16291_),
    .A2(_16297_),
    .B1(_16295_),
    .Y(_16348_));
 sky130_fd_sc_hd__nand3_4 _38925_ (.A(_16338_),
    .B(_16341_),
    .C(_16340_),
    .Y(_16349_));
 sky130_fd_sc_hd__nand3_2 _38926_ (.A(_16347_),
    .B(_16348_),
    .C(_16349_),
    .Y(_16350_));
 sky130_fd_sc_hd__nand3_4 _38927_ (.A(_16345_),
    .B(_16346_),
    .C(_16350_),
    .Y(_16351_));
 sky130_fd_sc_hd__o21ai_4 _38928_ (.A1(_16342_),
    .A2(_16344_),
    .B1(_16348_),
    .Y(_16352_));
 sky130_fd_sc_hd__a22oi_4 _38929_ (.A1(_16118_),
    .A2(_16132_),
    .B1(_16130_),
    .B2(_16134_),
    .Y(_16353_));
 sky130_fd_sc_hd__nand2_1 _38930_ (.A(_16291_),
    .B(_16293_),
    .Y(_16354_));
 sky130_fd_sc_hd__nand2_1 _38931_ (.A(_16354_),
    .B(_16296_),
    .Y(_16355_));
 sky130_fd_sc_hd__nand2_2 _38932_ (.A(_16355_),
    .B(_16298_),
    .Y(_16356_));
 sky130_fd_sc_hd__nand3_4 _38933_ (.A(_16347_),
    .B(_16356_),
    .C(_16349_),
    .Y(_16357_));
 sky130_fd_sc_hd__nand3_4 _38934_ (.A(_16352_),
    .B(_16353_),
    .C(_16357_),
    .Y(_16358_));
 sky130_fd_sc_hd__a21boi_4 _38935_ (.A1(_16066_),
    .A2(_16071_),
    .B1_N(_16070_),
    .Y(_16359_));
 sky130_fd_sc_hd__a31o_2 _38936_ (.A1(_20080_),
    .A2(_20084_),
    .A3(_16159_),
    .B1(_16058_),
    .X(_16360_));
 sky130_fd_sc_hd__nor2_8 _38937_ (.A(_16148_),
    .B(_16146_),
    .Y(_16361_));
 sky130_fd_sc_hd__o21a_2 _38938_ (.A1(_10067_),
    .A2(_07295_),
    .B1(net504),
    .X(_16362_));
 sky130_fd_sc_hd__nand2_2 _38939_ (.A(_16362_),
    .B(_06641_),
    .Y(_16363_));
 sky130_fd_sc_hd__or2_2 _38940_ (.A(_16361_),
    .B(_16363_),
    .X(_16364_));
 sky130_vsdinv _38941_ (.A(_16362_),
    .Y(_16365_));
 sky130_fd_sc_hd__o21ai_2 _38942_ (.A1(_16361_),
    .A2(_16365_),
    .B1(_15813_),
    .Y(_16366_));
 sky130_fd_sc_hd__and2_1 _38943_ (.A(_16364_),
    .B(_16366_),
    .X(_16367_));
 sky130_fd_sc_hd__clkbuf_4 _38944_ (.A(_16367_),
    .X(_16368_));
 sky130_fd_sc_hd__nor2_4 _38945_ (.A(_16360_),
    .B(_16368_),
    .Y(_16369_));
 sky130_vsdinv _38946_ (.A(_16369_),
    .Y(_16370_));
 sky130_fd_sc_hd__nand2_2 _38947_ (.A(_16152_),
    .B(_16150_),
    .Y(_16371_));
 sky130_vsdinv _38948_ (.A(_16371_),
    .Y(_16372_));
 sky130_fd_sc_hd__nand2_2 _38949_ (.A(_16368_),
    .B(_16360_),
    .Y(_16373_));
 sky130_fd_sc_hd__nand3_2 _38950_ (.A(_16370_),
    .B(_16372_),
    .C(_16373_),
    .Y(_16374_));
 sky130_fd_sc_hd__and3_1 _38951_ (.A(_16360_),
    .B(_16366_),
    .C(_16364_),
    .X(_16375_));
 sky130_fd_sc_hd__o21ai_2 _38952_ (.A1(_16369_),
    .A2(_16375_),
    .B1(_16371_),
    .Y(_16376_));
 sky130_fd_sc_hd__a21oi_4 _38953_ (.A1(_16156_),
    .A2(_16155_),
    .B1(_16154_),
    .Y(_16377_));
 sky130_fd_sc_hd__nand3_4 _38954_ (.A(_16374_),
    .B(_16376_),
    .C(_16377_),
    .Y(_16378_));
 sky130_fd_sc_hd__nand3_2 _38955_ (.A(_16370_),
    .B(_16371_),
    .C(_16373_),
    .Y(_16379_));
 sky130_fd_sc_hd__o21ai_2 _38956_ (.A1(_16369_),
    .A2(_16375_),
    .B1(_16372_),
    .Y(_16380_));
 sky130_fd_sc_hd__a21o_1 _38957_ (.A1(_16156_),
    .A2(_16155_),
    .B1(_16154_),
    .X(_16381_));
 sky130_fd_sc_hd__nand3_4 _38958_ (.A(_16379_),
    .B(_16380_),
    .C(_16381_),
    .Y(_16382_));
 sky130_fd_sc_hd__nand2_1 _38959_ (.A(_16378_),
    .B(_16382_),
    .Y(_16383_));
 sky130_fd_sc_hd__nand2_1 _38960_ (.A(_16383_),
    .B(_16170_),
    .Y(_16384_));
 sky130_fd_sc_hd__nand3_2 _38961_ (.A(_16378_),
    .B(_16382_),
    .C(_16172_),
    .Y(_16385_));
 sky130_fd_sc_hd__nand3b_4 _38962_ (.A_N(_16359_),
    .B(_16384_),
    .C(_16385_),
    .Y(_16386_));
 sky130_fd_sc_hd__buf_2 _38963_ (.A(_15835_),
    .X(_16387_));
 sky130_fd_sc_hd__nand2_1 _38964_ (.A(_16383_),
    .B(_16387_),
    .Y(_16388_));
 sky130_fd_sc_hd__buf_4 _38965_ (.A(_15840_),
    .X(_16389_));
 sky130_fd_sc_hd__nand3_2 _38966_ (.A(_16378_),
    .B(_16382_),
    .C(_16389_),
    .Y(_16390_));
 sky130_fd_sc_hd__nand3_4 _38967_ (.A(_16388_),
    .B(_16359_),
    .C(_16390_),
    .Y(_16391_));
 sky130_vsdinv _38968_ (.A(_16164_),
    .Y(_16392_));
 sky130_fd_sc_hd__a21oi_4 _38969_ (.A1(_16172_),
    .A2(_16168_),
    .B1(_16392_),
    .Y(_16393_));
 sky130_vsdinv _38970_ (.A(_16393_),
    .Y(_16394_));
 sky130_fd_sc_hd__a21oi_4 _38971_ (.A1(_16386_),
    .A2(_16391_),
    .B1(_16394_),
    .Y(_16395_));
 sky130_fd_sc_hd__nand2_2 _38972_ (.A(_16386_),
    .B(_16391_),
    .Y(_16396_));
 sky130_fd_sc_hd__nor2_4 _38973_ (.A(_16393_),
    .B(_16396_),
    .Y(_16397_));
 sky130_fd_sc_hd__o2bb2ai_4 _38974_ (.A1_N(_16351_),
    .A2_N(_16358_),
    .B1(_16395_),
    .B2(_16397_),
    .Y(_16398_));
 sky130_fd_sc_hd__nor2_2 _38975_ (.A(_16395_),
    .B(_16397_),
    .Y(_16399_));
 sky130_fd_sc_hd__nand3_4 _38976_ (.A(_16399_),
    .B(_16358_),
    .C(_16351_),
    .Y(_16400_));
 sky130_fd_sc_hd__nand2_4 _38977_ (.A(_16190_),
    .B(_16136_),
    .Y(_16401_));
 sky130_fd_sc_hd__a21oi_4 _38978_ (.A1(_16398_),
    .A2(_16400_),
    .B1(_16401_),
    .Y(_16402_));
 sky130_vsdinv _38979_ (.A(_16174_),
    .Y(_16403_));
 sky130_fd_sc_hd__nand2_1 _38980_ (.A(_16182_),
    .B(_16179_),
    .Y(_16404_));
 sky130_fd_sc_hd__o21ai_1 _38981_ (.A1(_16251_),
    .A2(_16403_),
    .B1(_16404_),
    .Y(_16405_));
 sky130_fd_sc_hd__a31oi_2 _38982_ (.A1(_16137_),
    .A2(_16141_),
    .A3(_16142_),
    .B1(_16405_),
    .Y(_16406_));
 sky130_fd_sc_hd__o211a_1 _38983_ (.A1(_16189_),
    .A2(_16406_),
    .B1(_16400_),
    .C1(_16398_),
    .X(_16407_));
 sky130_fd_sc_hd__o22ai_4 _38984_ (.A1(_16265_),
    .A2(_16267_),
    .B1(_16402_),
    .B2(_16407_),
    .Y(_16408_));
 sky130_fd_sc_hd__a21o_1 _38985_ (.A1(_16398_),
    .A2(_16400_),
    .B1(_16401_),
    .X(_16409_));
 sky130_fd_sc_hd__nand3_4 _38986_ (.A(_16401_),
    .B(_16398_),
    .C(_16400_),
    .Y(_16410_));
 sky130_fd_sc_hd__nor2_4 _38987_ (.A(_16267_),
    .B(_16265_),
    .Y(_16411_));
 sky130_fd_sc_hd__nand3_4 _38988_ (.A(_16409_),
    .B(_16410_),
    .C(_16411_),
    .Y(_16412_));
 sky130_fd_sc_hd__a22oi_4 _38989_ (.A1(_16196_),
    .A2(_16250_),
    .B1(_16408_),
    .B2(_16412_),
    .Y(_16413_));
 sky130_fd_sc_hd__a21oi_1 _38990_ (.A1(_16194_),
    .A2(_16195_),
    .B1(_16193_),
    .Y(_16414_));
 sky130_fd_sc_hd__o211a_2 _38991_ (.A1(_16191_),
    .A2(_16414_),
    .B1(_16412_),
    .C1(_16408_),
    .X(_16415_));
 sky130_fd_sc_hd__o22ai_4 _38992_ (.A1(_16248_),
    .A2(_16249_),
    .B1(_16413_),
    .B2(_16415_),
    .Y(_16416_));
 sky130_fd_sc_hd__o21ai_2 _38993_ (.A1(_16193_),
    .A2(_16188_),
    .B1(_16197_),
    .Y(_16417_));
 sky130_fd_sc_hd__a21o_2 _38994_ (.A1(_16408_),
    .A2(_16412_),
    .B1(_16417_),
    .X(_16418_));
 sky130_fd_sc_hd__nand3_4 _38995_ (.A(_16408_),
    .B(_16417_),
    .C(_16412_),
    .Y(_16419_));
 sky130_fd_sc_hd__nor2_4 _38996_ (.A(_16249_),
    .B(_16248_),
    .Y(_16420_));
 sky130_fd_sc_hd__nand3_2 _38997_ (.A(_16418_),
    .B(_16419_),
    .C(_16420_),
    .Y(_16421_));
 sky130_fd_sc_hd__nand3_4 _38998_ (.A(_16246_),
    .B(_16416_),
    .C(_16421_),
    .Y(_16422_));
 sky130_fd_sc_hd__buf_6 _38999_ (.A(_14930_),
    .X(_16423_));
 sky130_fd_sc_hd__nand2_4 _39000_ (.A(_16247_),
    .B(_16423_),
    .Y(_16424_));
 sky130_vsdinv _39001_ (.A(_16424_),
    .Y(_16425_));
 sky130_fd_sc_hd__buf_4 _39002_ (.A(_14931_),
    .X(_16426_));
 sky130_fd_sc_hd__nor2_2 _39003_ (.A(_16426_),
    .B(_16247_),
    .Y(_16427_));
 sky130_fd_sc_hd__o22ai_4 _39004_ (.A1(_16425_),
    .A2(_16427_),
    .B1(_16413_),
    .B2(_16415_),
    .Y(_16428_));
 sky130_fd_sc_hd__o21ai_2 _39005_ (.A1(_16208_),
    .A2(_16201_),
    .B1(_16213_),
    .Y(_16429_));
 sky130_vsdinv _39006_ (.A(_16420_),
    .Y(_16430_));
 sky130_fd_sc_hd__nand3_4 _39007_ (.A(_16418_),
    .B(_16419_),
    .C(_16430_),
    .Y(_16431_));
 sky130_fd_sc_hd__nand3_4 _39008_ (.A(_16428_),
    .B(_16429_),
    .C(_16431_),
    .Y(_16432_));
 sky130_fd_sc_hd__nand2_1 _39009_ (.A(_16422_),
    .B(_16432_),
    .Y(_16433_));
 sky130_fd_sc_hd__nand2_1 _39010_ (.A(_16433_),
    .B(_16205_),
    .Y(_16434_));
 sky130_fd_sc_hd__nand3_2 _39011_ (.A(_16422_),
    .B(_16432_),
    .C(_16206_),
    .Y(_16435_));
 sky130_fd_sc_hd__nand3_4 _39012_ (.A(_16245_),
    .B(_16434_),
    .C(_16435_),
    .Y(_16436_));
 sky130_fd_sc_hd__nand3_4 _39013_ (.A(_16422_),
    .B(_16432_),
    .C(_16205_),
    .Y(_16437_));
 sky130_fd_sc_hd__nand2_1 _39014_ (.A(_16433_),
    .B(_16206_),
    .Y(_16438_));
 sky130_fd_sc_hd__o211ai_4 _39015_ (.A1(_16225_),
    .A2(_16244_),
    .B1(_16437_),
    .C1(_16438_),
    .Y(_16439_));
 sky130_fd_sc_hd__and2_1 _39016_ (.A(_16436_),
    .B(_16439_),
    .X(_16440_));
 sky130_fd_sc_hd__a21bo_1 _39017_ (.A1(_16242_),
    .A2(_16224_),
    .B1_N(_16228_),
    .X(_16441_));
 sky130_fd_sc_hd__xor2_1 _39018_ (.A(_16440_),
    .B(_16441_),
    .X(_02668_));
 sky130_fd_sc_hd__o21ai_2 _39019_ (.A1(_16342_),
    .A2(_16356_),
    .B1(_16349_),
    .Y(_16442_));
 sky130_fd_sc_hd__a21oi_4 _39020_ (.A1(_16315_),
    .A2(_16316_),
    .B1(_16300_),
    .Y(_16443_));
 sky130_fd_sc_hd__nand2_1 _39021_ (.A(_16336_),
    .B(_16332_),
    .Y(_16444_));
 sky130_fd_sc_hd__a31oi_4 _39022_ (.A1(_16315_),
    .A2(_16300_),
    .A3(_16316_),
    .B1(_16444_),
    .Y(_16445_));
 sky130_fd_sc_hd__nor2_4 _39023_ (.A(net441),
    .B(_15929_),
    .Y(_16446_));
 sky130_fd_sc_hd__and4_2 _39024_ (.A(_10691_),
    .B(_13837_),
    .C(_19830_),
    .D(_20115_),
    .X(_16447_));
 sky130_fd_sc_hd__clkbuf_2 _39025_ (.A(_13142_),
    .X(_16448_));
 sky130_fd_sc_hd__o22a_2 _39026_ (.A1(_20120_),
    .A2(_16448_),
    .B1(_16102_),
    .B2(_11074_),
    .X(_16449_));
 sky130_fd_sc_hd__or3_4 _39027_ (.A(_16446_),
    .B(_16447_),
    .C(_16449_),
    .X(_16450_));
 sky130_fd_sc_hd__o21ai_4 _39028_ (.A1(_16447_),
    .A2(_16449_),
    .B1(_16446_),
    .Y(_16451_));
 sky130_fd_sc_hd__o21ba_2 _39029_ (.A1(_16304_),
    .A2(_16302_),
    .B1_N(_16301_),
    .X(_16452_));
 sky130_fd_sc_hd__a21oi_1 _39030_ (.A1(_16450_),
    .A2(_16451_),
    .B1(_16452_),
    .Y(_16453_));
 sky130_fd_sc_hd__and3_1 _39031_ (.A(_16450_),
    .B(_16451_),
    .C(_16452_),
    .X(_16454_));
 sky130_fd_sc_hd__o22a_2 _39032_ (.A1(_16094_),
    .A2(_09733_),
    .B1(_16095_),
    .B2(_12100_),
    .X(_16455_));
 sky130_fd_sc_hd__a31o_1 _39033_ (.A1(_20106_),
    .A2(_20109_),
    .A3(_16093_),
    .B1(_16455_),
    .X(_16456_));
 sky130_fd_sc_hd__nand2_2 _39034_ (.A(_15897_),
    .B(_20103_),
    .Y(_16457_));
 sky130_vsdinv _39035_ (.A(_16457_),
    .Y(_16458_));
 sky130_fd_sc_hd__nand2_1 _39036_ (.A(_16456_),
    .B(_16458_),
    .Y(_16459_));
 sky130_fd_sc_hd__and3_1 _39037_ (.A(_16092_),
    .B(_20106_),
    .C(_13758_),
    .X(_16460_));
 sky130_fd_sc_hd__nor2_1 _39038_ (.A(_16455_),
    .B(_16460_),
    .Y(_16461_));
 sky130_fd_sc_hd__nand2_1 _39039_ (.A(_16461_),
    .B(_16457_),
    .Y(_16462_));
 sky130_fd_sc_hd__nand2_2 _39040_ (.A(_16459_),
    .B(_16462_),
    .Y(_16463_));
 sky130_fd_sc_hd__o21ai_2 _39041_ (.A1(_16453_),
    .A2(_16454_),
    .B1(_16463_),
    .Y(_16464_));
 sky130_vsdinv _39042_ (.A(_16463_),
    .Y(_16465_));
 sky130_fd_sc_hd__a21o_1 _39043_ (.A1(_16450_),
    .A2(_16451_),
    .B1(_16452_),
    .X(_16466_));
 sky130_fd_sc_hd__nand3_4 _39044_ (.A(_16450_),
    .B(_16451_),
    .C(_16452_),
    .Y(_16467_));
 sky130_fd_sc_hd__nand3_4 _39045_ (.A(_16465_),
    .B(_16466_),
    .C(_16467_),
    .Y(_16468_));
 sky130_vsdinv _39046_ (.A(_16314_),
    .Y(_16469_));
 sky130_fd_sc_hd__a21oi_2 _39047_ (.A1(_16303_),
    .A2(_16305_),
    .B1(_16306_),
    .Y(_16470_));
 sky130_fd_sc_hd__a21oi_4 _39048_ (.A1(_16469_),
    .A2(_16308_),
    .B1(_16470_),
    .Y(_16471_));
 sky130_fd_sc_hd__a21o_4 _39049_ (.A1(_16464_),
    .A2(_16468_),
    .B1(_16471_),
    .X(_16472_));
 sky130_fd_sc_hd__nand2_1 _39050_ (.A(_19855_),
    .B(_20092_),
    .Y(_16473_));
 sky130_fd_sc_hd__nand2_1 _39051_ (.A(_15597_),
    .B(_20098_),
    .Y(_16474_));
 sky130_fd_sc_hd__nand2_1 _39052_ (.A(_15594_),
    .B(_13451_),
    .Y(_16475_));
 sky130_fd_sc_hd__nor2_1 _39053_ (.A(_16474_),
    .B(_16475_),
    .Y(_16476_));
 sky130_fd_sc_hd__nand2_1 _39054_ (.A(_16474_),
    .B(_16475_),
    .Y(_16477_));
 sky130_fd_sc_hd__or3b_4 _39055_ (.A(_16473_),
    .B(_16476_),
    .C_N(_16477_),
    .X(_16478_));
 sky130_vsdinv _39056_ (.A(_16476_),
    .Y(_16479_));
 sky130_fd_sc_hd__a21bo_1 _39057_ (.A1(_16479_),
    .A2(_16477_),
    .B1_N(_16473_),
    .X(_16480_));
 sky130_fd_sc_hd__a32o_2 _39058_ (.A1(_16093_),
    .A2(_20109_),
    .A3(_20112_),
    .B1(_16312_),
    .B2(_16310_),
    .X(_16481_));
 sky130_fd_sc_hd__a21o_1 _39059_ (.A1(_16478_),
    .A2(_16480_),
    .B1(_16481_),
    .X(_16482_));
 sky130_fd_sc_hd__nand3_4 _39060_ (.A(_16478_),
    .B(_16481_),
    .C(_16480_),
    .Y(_16483_));
 sky130_vsdinv _39061_ (.A(_16326_),
    .Y(_16484_));
 sky130_fd_sc_hd__nor2_2 _39062_ (.A(_16322_),
    .B(_16484_),
    .Y(_16485_));
 sky130_fd_sc_hd__a21boi_4 _39063_ (.A1(_16482_),
    .A2(_16483_),
    .B1_N(_16485_),
    .Y(_16486_));
 sky130_fd_sc_hd__o211a_2 _39064_ (.A1(_16322_),
    .A2(_16484_),
    .B1(_16483_),
    .C1(_16482_),
    .X(_16487_));
 sky130_fd_sc_hd__nor2_4 _39065_ (.A(_16486_),
    .B(_16487_),
    .Y(_16488_));
 sky130_fd_sc_hd__nand3_4 _39066_ (.A(_16464_),
    .B(_16471_),
    .C(_16468_),
    .Y(_16489_));
 sky130_fd_sc_hd__nand3_4 _39067_ (.A(_16472_),
    .B(_16488_),
    .C(_16489_),
    .Y(_16490_));
 sky130_fd_sc_hd__o2bb2ai_2 _39068_ (.A1_N(_16489_),
    .A2_N(_16472_),
    .B1(_16486_),
    .B2(_16487_),
    .Y(_16491_));
 sky130_fd_sc_hd__o211ai_4 _39069_ (.A1(_16443_),
    .A2(_16445_),
    .B1(_16490_),
    .C1(_16491_),
    .Y(_16492_));
 sky130_fd_sc_hd__nand2_1 _39070_ (.A(_16472_),
    .B(_16489_),
    .Y(_16493_));
 sky130_fd_sc_hd__nand2_1 _39071_ (.A(_16493_),
    .B(_16488_),
    .Y(_16494_));
 sky130_fd_sc_hd__a21oi_4 _39072_ (.A1(_16339_),
    .A2(_16317_),
    .B1(_16443_),
    .Y(_16495_));
 sky130_fd_sc_hd__nand3b_2 _39073_ (.A_N(_16488_),
    .B(_16472_),
    .C(_16489_),
    .Y(_16496_));
 sky130_fd_sc_hd__nand3_4 _39074_ (.A(_16494_),
    .B(_16495_),
    .C(_16496_),
    .Y(_16497_));
 sky130_fd_sc_hd__nand2_2 _39075_ (.A(_19867_),
    .B(_13647_),
    .Y(_16498_));
 sky130_fd_sc_hd__nand2_1 _39076_ (.A(_11396_),
    .B(_20087_),
    .Y(_16499_));
 sky130_fd_sc_hd__nand2_1 _39077_ (.A(_12855_),
    .B(_12298_),
    .Y(_16500_));
 sky130_fd_sc_hd__nor2_2 _39078_ (.A(_16499_),
    .B(_16500_),
    .Y(_16501_));
 sky130_fd_sc_hd__and2_1 _39079_ (.A(_16499_),
    .B(_16500_),
    .X(_16502_));
 sky130_fd_sc_hd__or3_4 _39080_ (.A(_16498_),
    .B(_16501_),
    .C(_16502_),
    .X(_16503_));
 sky130_fd_sc_hd__o21ai_2 _39081_ (.A1(_16501_),
    .A2(_16502_),
    .B1(_16498_),
    .Y(_16504_));
 sky130_fd_sc_hd__nand2_2 _39082_ (.A(_16276_),
    .B(_16272_),
    .Y(_16505_));
 sky130_fd_sc_hd__a21oi_1 _39083_ (.A1(_16503_),
    .A2(_16504_),
    .B1(_16505_),
    .Y(_16506_));
 sky130_fd_sc_hd__nand3_4 _39084_ (.A(_16503_),
    .B(_16504_),
    .C(_16505_),
    .Y(_16507_));
 sky130_vsdinv _39085_ (.A(_16507_),
    .Y(_16508_));
 sky130_fd_sc_hd__nand2_4 _39086_ (.A(_11603_),
    .B(net457),
    .Y(_16509_));
 sky130_vsdinv _39087_ (.A(_16509_),
    .Y(_16510_));
 sky130_fd_sc_hd__and4_1 _39088_ (.A(_19871_),
    .B(_10945_),
    .C(_11604_),
    .D(_20074_),
    .X(_16511_));
 sky130_vsdinv _39089_ (.A(_19871_),
    .Y(_16512_));
 sky130_fd_sc_hd__nand2_1 _39090_ (.A(_19875_),
    .B(_11604_),
    .Y(_16513_));
 sky130_fd_sc_hd__o21a_1 _39091_ (.A1(_16512_),
    .A2(_10767_),
    .B1(_16513_),
    .X(_16514_));
 sky130_fd_sc_hd__nor2_1 _39092_ (.A(_16511_),
    .B(_16514_),
    .Y(_16515_));
 sky130_fd_sc_hd__or2_1 _39093_ (.A(_16510_),
    .B(_16515_),
    .X(_16516_));
 sky130_fd_sc_hd__nand2_1 _39094_ (.A(_16515_),
    .B(_16510_),
    .Y(_16517_));
 sky130_fd_sc_hd__nand2_1 _39095_ (.A(_16516_),
    .B(_16517_),
    .Y(_16518_));
 sky130_fd_sc_hd__o21ai_2 _39096_ (.A1(_16506_),
    .A2(_16508_),
    .B1(_16518_),
    .Y(_16519_));
 sky130_fd_sc_hd__a21o_1 _39097_ (.A1(_16503_),
    .A2(_16504_),
    .B1(_16505_),
    .X(_16520_));
 sky130_fd_sc_hd__nand3b_4 _39098_ (.A_N(_16518_),
    .B(_16507_),
    .C(_16520_),
    .Y(_16521_));
 sky130_fd_sc_hd__nand2_1 _39099_ (.A(_16519_),
    .B(_16521_),
    .Y(_16522_));
 sky130_fd_sc_hd__a21boi_1 _39100_ (.A1(_16329_),
    .A2(_16330_),
    .B1_N(_16331_),
    .Y(_16523_));
 sky130_fd_sc_hd__nand2_2 _39101_ (.A(_16522_),
    .B(_16523_),
    .Y(_16524_));
 sky130_fd_sc_hd__nand2_1 _39102_ (.A(_16332_),
    .B(_16331_),
    .Y(_16525_));
 sky130_fd_sc_hd__nand3_4 _39103_ (.A(_16525_),
    .B(_16519_),
    .C(_16521_),
    .Y(_16526_));
 sky130_vsdinv _39104_ (.A(_16286_),
    .Y(_16527_));
 sky130_fd_sc_hd__a21bo_1 _39105_ (.A1(_16278_),
    .A2(_16527_),
    .B1_N(_16279_),
    .X(_16528_));
 sky130_fd_sc_hd__and3_2 _39106_ (.A(_16524_),
    .B(_16526_),
    .C(_16528_),
    .X(_16529_));
 sky130_fd_sc_hd__a21oi_4 _39107_ (.A1(_16524_),
    .A2(_16526_),
    .B1(_16528_),
    .Y(_16530_));
 sky130_fd_sc_hd__o2bb2ai_2 _39108_ (.A1_N(_16492_),
    .A2_N(_16497_),
    .B1(_16529_),
    .B2(_16530_),
    .Y(_16531_));
 sky130_fd_sc_hd__nor2_8 _39109_ (.A(_16530_),
    .B(_16529_),
    .Y(_16532_));
 sky130_fd_sc_hd__nand3_4 _39110_ (.A(_16497_),
    .B(_16492_),
    .C(_16532_),
    .Y(_16533_));
 sky130_fd_sc_hd__nand3_4 _39111_ (.A(_16442_),
    .B(_16531_),
    .C(_16533_),
    .Y(_16534_));
 sky130_fd_sc_hd__a21oi_4 _39112_ (.A1(_16347_),
    .A2(_16348_),
    .B1(_16344_),
    .Y(_16535_));
 sky130_fd_sc_hd__nand2_1 _39113_ (.A(_16497_),
    .B(_16492_),
    .Y(_16536_));
 sky130_fd_sc_hd__nand2_1 _39114_ (.A(_16536_),
    .B(_16532_),
    .Y(_16537_));
 sky130_fd_sc_hd__nand3b_2 _39115_ (.A_N(_16532_),
    .B(_16497_),
    .C(_16492_),
    .Y(_16538_));
 sky130_fd_sc_hd__nand3_4 _39116_ (.A(_16535_),
    .B(_16537_),
    .C(_16538_),
    .Y(_16539_));
 sky130_fd_sc_hd__a21oi_4 _39117_ (.A1(_16292_),
    .A2(_16288_),
    .B1(_16290_),
    .Y(_16540_));
 sky130_fd_sc_hd__a31o_2 _39118_ (.A1(_20075_),
    .A2(_20080_),
    .A3(_16159_),
    .B1(_16284_),
    .X(_16541_));
 sky130_fd_sc_hd__or2_2 _39119_ (.A(_16541_),
    .B(_16368_),
    .X(_16542_));
 sky130_fd_sc_hd__nand2_2 _39120_ (.A(_16368_),
    .B(_16541_),
    .Y(_16543_));
 sky130_vsdinv _39121_ (.A(_16361_),
    .Y(_16544_));
 sky130_fd_sc_hd__nand2_4 _39122_ (.A(_16544_),
    .B(_16363_),
    .Y(_16545_));
 sky130_fd_sc_hd__nand3_2 _39123_ (.A(_16542_),
    .B(_16543_),
    .C(_16545_),
    .Y(_16546_));
 sky130_fd_sc_hd__nor2_4 _39124_ (.A(_16541_),
    .B(_16368_),
    .Y(_16547_));
 sky130_fd_sc_hd__and3_1 _39125_ (.A(_16541_),
    .B(_16366_),
    .C(_16364_),
    .X(_16548_));
 sky130_vsdinv _39126_ (.A(_16545_),
    .Y(_16549_));
 sky130_fd_sc_hd__o21ai_2 _39127_ (.A1(_16547_),
    .A2(_16548_),
    .B1(_16549_),
    .Y(_16550_));
 sky130_fd_sc_hd__o21ai_2 _39128_ (.A1(_16372_),
    .A2(_16369_),
    .B1(_16373_),
    .Y(_16551_));
 sky130_fd_sc_hd__nand3_4 _39129_ (.A(_16546_),
    .B(_16550_),
    .C(_16551_),
    .Y(_16552_));
 sky130_vsdinv _39130_ (.A(_16552_),
    .Y(_16553_));
 sky130_fd_sc_hd__nand3_2 _39131_ (.A(_16542_),
    .B(_16543_),
    .C(_16549_),
    .Y(_16554_));
 sky130_fd_sc_hd__o21ai_2 _39132_ (.A1(_16547_),
    .A2(_16548_),
    .B1(_16545_),
    .Y(_16555_));
 sky130_fd_sc_hd__nand3b_4 _39133_ (.A_N(_16551_),
    .B(_16554_),
    .C(_16555_),
    .Y(_16556_));
 sky130_fd_sc_hd__nand2_2 _39134_ (.A(_16556_),
    .B(_16172_),
    .Y(_16557_));
 sky130_fd_sc_hd__nand2_1 _39135_ (.A(_16556_),
    .B(_16552_),
    .Y(_16558_));
 sky130_fd_sc_hd__nand2_1 _39136_ (.A(_16558_),
    .B(_16389_),
    .Y(_16559_));
 sky130_fd_sc_hd__o221ai_4 _39137_ (.A1(_16540_),
    .A2(_16297_),
    .B1(_16553_),
    .B2(_16557_),
    .C1(_16559_),
    .Y(_16560_));
 sky130_fd_sc_hd__nor2_4 _39138_ (.A(_16540_),
    .B(_16297_),
    .Y(_16561_));
 sky130_fd_sc_hd__nand2_2 _39139_ (.A(_16558_),
    .B(_16387_),
    .Y(_16562_));
 sky130_fd_sc_hd__nand3_4 _39140_ (.A(_16556_),
    .B(_16552_),
    .C(_16389_),
    .Y(_16563_));
 sky130_fd_sc_hd__nand3_4 _39141_ (.A(_16561_),
    .B(_16562_),
    .C(_16563_),
    .Y(_16564_));
 sky130_vsdinv _39142_ (.A(_16382_),
    .Y(_16565_));
 sky130_fd_sc_hd__a21o_1 _39143_ (.A1(_16387_),
    .A2(_16378_),
    .B1(_16565_),
    .X(_16566_));
 sky130_fd_sc_hd__a21oi_4 _39144_ (.A1(_16560_),
    .A2(_16564_),
    .B1(_16566_),
    .Y(_16567_));
 sky130_fd_sc_hd__nand3_4 _39145_ (.A(_16560_),
    .B(_16564_),
    .C(_16566_),
    .Y(_16568_));
 sky130_vsdinv _39146_ (.A(_16568_),
    .Y(_16569_));
 sky130_fd_sc_hd__o2bb2ai_4 _39147_ (.A1_N(_16534_),
    .A2_N(_16539_),
    .B1(_16567_),
    .B2(_16569_),
    .Y(_16570_));
 sky130_fd_sc_hd__a21oi_2 _39148_ (.A1(_16387_),
    .A2(_16378_),
    .B1(_16565_),
    .Y(_16571_));
 sky130_fd_sc_hd__a21oi_4 _39149_ (.A1(_16562_),
    .A2(_16563_),
    .B1(_16561_),
    .Y(_16572_));
 sky130_fd_sc_hd__nor2_2 _39150_ (.A(_16571_),
    .B(_16572_),
    .Y(_16573_));
 sky130_fd_sc_hd__a21oi_4 _39151_ (.A1(_16573_),
    .A2(_16564_),
    .B1(_16567_),
    .Y(_16574_));
 sky130_fd_sc_hd__nand3_4 _39152_ (.A(_16539_),
    .B(_16534_),
    .C(_16574_),
    .Y(_16575_));
 sky130_fd_sc_hd__nand2_1 _39153_ (.A(_16399_),
    .B(_16358_),
    .Y(_16576_));
 sky130_fd_sc_hd__nand2_2 _39154_ (.A(_16576_),
    .B(_16351_),
    .Y(_16577_));
 sky130_fd_sc_hd__a21oi_4 _39155_ (.A1(_16570_),
    .A2(_16575_),
    .B1(_16577_),
    .Y(_16578_));
 sky130_vsdinv _39156_ (.A(_16351_),
    .Y(_16579_));
 sky130_fd_sc_hd__nand2_1 _39157_ (.A(_16396_),
    .B(_16393_),
    .Y(_16580_));
 sky130_fd_sc_hd__nand3_2 _39158_ (.A(_16386_),
    .B(_16394_),
    .C(_16391_),
    .Y(_16581_));
 sky130_fd_sc_hd__nand2_1 _39159_ (.A(_16580_),
    .B(_16581_),
    .Y(_16582_));
 sky130_fd_sc_hd__a31oi_4 _39160_ (.A1(_16353_),
    .A2(_16352_),
    .A3(_16357_),
    .B1(_16582_),
    .Y(_16583_));
 sky130_fd_sc_hd__o211a_2 _39161_ (.A1(_16579_),
    .A2(_16583_),
    .B1(_16575_),
    .C1(_16570_),
    .X(_16584_));
 sky130_fd_sc_hd__nand3_2 _39162_ (.A(_16581_),
    .B(_16386_),
    .C(_16258_),
    .Y(_16585_));
 sky130_fd_sc_hd__nor2_1 _39163_ (.A(_14009_),
    .B(_16252_),
    .Y(_16586_));
 sky130_fd_sc_hd__or2_4 _39164_ (.A(_16253_),
    .B(_16586_),
    .X(_16587_));
 sky130_vsdinv _39165_ (.A(_16587_),
    .Y(_16588_));
 sky130_fd_sc_hd__nand2_1 _39166_ (.A(_16585_),
    .B(_16588_),
    .Y(_16589_));
 sky130_fd_sc_hd__a21o_1 _39167_ (.A1(_16581_),
    .A2(_16386_),
    .B1(_16258_),
    .X(_16590_));
 sky130_fd_sc_hd__or2b_2 _39168_ (.A(_16589_),
    .B_N(_16590_),
    .X(_16591_));
 sky130_fd_sc_hd__clkbuf_4 _39169_ (.A(_16588_),
    .X(_16592_));
 sky130_fd_sc_hd__a21o_1 _39170_ (.A1(_16590_),
    .A2(_16585_),
    .B1(_16592_),
    .X(_16593_));
 sky130_fd_sc_hd__nand2_4 _39171_ (.A(_16591_),
    .B(_16593_),
    .Y(_16594_));
 sky130_fd_sc_hd__o21ai_2 _39172_ (.A1(_16578_),
    .A2(_16584_),
    .B1(_16594_),
    .Y(_16595_));
 sky130_fd_sc_hd__or2b_1 _39173_ (.A(_16267_),
    .B_N(_16264_),
    .X(_16596_));
 sky130_fd_sc_hd__o21ai_2 _39174_ (.A1(_16596_),
    .A2(_16402_),
    .B1(_16410_),
    .Y(_16597_));
 sky130_fd_sc_hd__nand2_1 _39175_ (.A(_16570_),
    .B(_16575_),
    .Y(_16598_));
 sky130_fd_sc_hd__nor2_2 _39176_ (.A(_16579_),
    .B(_16583_),
    .Y(_16599_));
 sky130_fd_sc_hd__nand2_2 _39177_ (.A(_16598_),
    .B(_16599_),
    .Y(_16600_));
 sky130_fd_sc_hd__and2_1 _39178_ (.A(_16591_),
    .B(_16593_),
    .X(_16601_));
 sky130_fd_sc_hd__nand3_4 _39179_ (.A(_16577_),
    .B(_16570_),
    .C(_16575_),
    .Y(_16602_));
 sky130_fd_sc_hd__nand3_2 _39180_ (.A(_16600_),
    .B(_16601_),
    .C(_16602_),
    .Y(_16603_));
 sky130_fd_sc_hd__nand3_4 _39181_ (.A(_16595_),
    .B(_16597_),
    .C(_16603_),
    .Y(_16604_));
 sky130_fd_sc_hd__o21ai_4 _39182_ (.A1(_16578_),
    .A2(_16584_),
    .B1(_16601_),
    .Y(_16605_));
 sky130_fd_sc_hd__a21oi_2 _39183_ (.A1(_16409_),
    .A2(_16411_),
    .B1(_16407_),
    .Y(_16606_));
 sky130_fd_sc_hd__nand3_4 _39184_ (.A(_16600_),
    .B(_16594_),
    .C(_16602_),
    .Y(_16607_));
 sky130_fd_sc_hd__nand3_4 _39185_ (.A(_16605_),
    .B(_16606_),
    .C(_16607_),
    .Y(_16608_));
 sky130_fd_sc_hd__nand2_1 _39186_ (.A(_16266_),
    .B(_16260_),
    .Y(_16609_));
 sky130_fd_sc_hd__nand2_2 _39187_ (.A(_16609_),
    .B(_16259_),
    .Y(_16610_));
 sky130_fd_sc_hd__nor2_2 _39188_ (.A(_15754_),
    .B(_16610_),
    .Y(_16611_));
 sky130_vsdinv _39189_ (.A(_16610_),
    .Y(_16612_));
 sky130_fd_sc_hd__nor2_2 _39190_ (.A(_14931_),
    .B(_16612_),
    .Y(_16613_));
 sky130_fd_sc_hd__o2bb2ai_4 _39191_ (.A1_N(_16604_),
    .A2_N(_16608_),
    .B1(_16611_),
    .B2(_16613_),
    .Y(_16614_));
 sky130_fd_sc_hd__or2_2 _39192_ (.A(_16611_),
    .B(_16613_),
    .X(_16615_));
 sky130_fd_sc_hd__nand3b_4 _39193_ (.A_N(_16615_),
    .B(_16608_),
    .C(_16604_),
    .Y(_16616_));
 sky130_fd_sc_hd__nand2_1 _39194_ (.A(_16419_),
    .B(_16420_),
    .Y(_16617_));
 sky130_fd_sc_hd__nand2_4 _39195_ (.A(_16617_),
    .B(_16418_),
    .Y(_16618_));
 sky130_fd_sc_hd__a21oi_4 _39196_ (.A1(_16614_),
    .A2(_16616_),
    .B1(_16618_),
    .Y(_16619_));
 sky130_fd_sc_hd__nand3_4 _39197_ (.A(_16614_),
    .B(_16618_),
    .C(_16616_),
    .Y(_16620_));
 sky130_fd_sc_hd__nand2_1 _39198_ (.A(_16620_),
    .B(_16425_),
    .Y(_16621_));
 sky130_vsdinv _39199_ (.A(_16428_),
    .Y(_16622_));
 sky130_fd_sc_hd__nand2_1 _39200_ (.A(_16429_),
    .B(_16431_),
    .Y(_16623_));
 sky130_fd_sc_hd__o2bb2ai_2 _39201_ (.A1_N(_16205_),
    .A2_N(_16422_),
    .B1(_16622_),
    .B2(_16623_),
    .Y(_16624_));
 sky130_fd_sc_hd__a21o_1 _39202_ (.A1(_16608_),
    .A2(_16604_),
    .B1(_16615_),
    .X(_16625_));
 sky130_fd_sc_hd__o21ai_2 _39203_ (.A1(_16420_),
    .A2(_16413_),
    .B1(_16419_),
    .Y(_16626_));
 sky130_fd_sc_hd__nand3_2 _39204_ (.A(_16608_),
    .B(_16604_),
    .C(_16615_),
    .Y(_16627_));
 sky130_fd_sc_hd__nand3_4 _39205_ (.A(_16625_),
    .B(_16626_),
    .C(_16627_),
    .Y(_16628_));
 sky130_fd_sc_hd__nand2_1 _39206_ (.A(_16628_),
    .B(_16620_),
    .Y(_16629_));
 sky130_fd_sc_hd__nand2_1 _39207_ (.A(_16629_),
    .B(_16424_),
    .Y(_16630_));
 sky130_fd_sc_hd__o211ai_4 _39208_ (.A1(_16619_),
    .A2(_16621_),
    .B1(_16624_),
    .C1(_16630_),
    .Y(_16631_));
 sky130_fd_sc_hd__nand2_2 _39209_ (.A(_16629_),
    .B(_16425_),
    .Y(_16632_));
 sky130_fd_sc_hd__a21boi_2 _39210_ (.A1(_16422_),
    .A2(_16205_),
    .B1_N(_16432_),
    .Y(_16633_));
 sky130_fd_sc_hd__nand3_4 _39211_ (.A(_16628_),
    .B(_16620_),
    .C(_16424_),
    .Y(_16634_));
 sky130_fd_sc_hd__nand3_4 _39212_ (.A(_16632_),
    .B(_16633_),
    .C(_16634_),
    .Y(_16635_));
 sky130_fd_sc_hd__nand2_1 _39213_ (.A(_16631_),
    .B(_16635_),
    .Y(_16636_));
 sky130_vsdinv _39214_ (.A(_16437_),
    .Y(_16637_));
 sky130_fd_sc_hd__o2bb2ai_2 _39215_ (.A1_N(_16206_),
    .A2_N(_16433_),
    .B1(_16225_),
    .B2(_16244_),
    .Y(_16638_));
 sky130_fd_sc_hd__o2111ai_4 _39216_ (.A1(_16637_),
    .A2(_16638_),
    .B1(_16228_),
    .C1(_16436_),
    .D1(_16224_),
    .Y(_16639_));
 sky130_vsdinv _39217_ (.A(_16639_),
    .Y(_16640_));
 sky130_fd_sc_hd__a21boi_4 _39218_ (.A1(_16228_),
    .A2(_16439_),
    .B1_N(_16436_),
    .Y(_16641_));
 sky130_fd_sc_hd__a21oi_2 _39219_ (.A1(_16242_),
    .A2(_16640_),
    .B1(_16641_),
    .Y(_16642_));
 sky130_fd_sc_hd__xor2_1 _39220_ (.A(_16636_),
    .B(_16642_),
    .X(_02669_));
 sky130_fd_sc_hd__a21oi_2 _39221_ (.A1(_16598_),
    .A2(_16599_),
    .B1(_16594_),
    .Y(_16643_));
 sky130_fd_sc_hd__nor2_4 _39222_ (.A(_10405_),
    .B(_12093_),
    .Y(_16644_));
 sky130_fd_sc_hd__and4_2 _39223_ (.A(_11074_),
    .B(_18695_),
    .C(_19830_),
    .D(_11492_),
    .X(_16645_));
 sky130_fd_sc_hd__o22a_2 _39224_ (.A1(_20115_),
    .A2(_16448_),
    .B1(_15916_),
    .B2(_15929_),
    .X(_16646_));
 sky130_fd_sc_hd__or3_4 _39225_ (.A(_16644_),
    .B(_16645_),
    .C(_16646_),
    .X(_16647_));
 sky130_fd_sc_hd__o21ai_4 _39226_ (.A1(_16645_),
    .A2(_16646_),
    .B1(_16644_),
    .Y(_16648_));
 sky130_fd_sc_hd__nor2_1 _39227_ (.A(_16446_),
    .B(_16447_),
    .Y(_16649_));
 sky130_fd_sc_hd__or2_4 _39228_ (.A(_16449_),
    .B(_16649_),
    .X(_16650_));
 sky130_fd_sc_hd__a21o_1 _39229_ (.A1(_16647_),
    .A2(_16648_),
    .B1(_16650_),
    .X(_16651_));
 sky130_fd_sc_hd__nand3_4 _39230_ (.A(_16650_),
    .B(_16648_),
    .C(_16647_),
    .Y(_16652_));
 sky130_fd_sc_hd__nand2_1 _39231_ (.A(_16651_),
    .B(_16652_),
    .Y(_16653_));
 sky130_fd_sc_hd__nand2_1 _39232_ (.A(_19844_),
    .B(_20099_),
    .Y(_16654_));
 sky130_vsdinv _39233_ (.A(_16654_),
    .Y(_16655_));
 sky130_fd_sc_hd__a22o_1 _39234_ (.A1(_15924_),
    .A2(_20106_),
    .B1(_15925_),
    .B2(_12303_),
    .X(_16656_));
 sky130_fd_sc_hd__o31ai_4 _39235_ (.A1(_16311_),
    .A2(_12604_),
    .A3(_12100_),
    .B1(_16656_),
    .Y(_16657_));
 sky130_fd_sc_hd__xor2_4 _39236_ (.A(_16655_),
    .B(_16657_),
    .X(_16658_));
 sky130_fd_sc_hd__nand2_1 _39237_ (.A(_16653_),
    .B(_16658_),
    .Y(_16659_));
 sky130_fd_sc_hd__nand2_1 _39238_ (.A(_16467_),
    .B(_16463_),
    .Y(_16660_));
 sky130_fd_sc_hd__nand2_1 _39239_ (.A(_16660_),
    .B(_16466_),
    .Y(_16661_));
 sky130_vsdinv _39240_ (.A(_16658_),
    .Y(_16662_));
 sky130_fd_sc_hd__nand3_2 _39241_ (.A(_16651_),
    .B(_16652_),
    .C(_16662_),
    .Y(_16663_));
 sky130_fd_sc_hd__nand3_4 _39242_ (.A(_16659_),
    .B(_16661_),
    .C(_16663_),
    .Y(_16664_));
 sky130_fd_sc_hd__nand2_2 _39243_ (.A(_16653_),
    .B(_16662_),
    .Y(_16665_));
 sky130_fd_sc_hd__and2_2 _39244_ (.A(_16660_),
    .B(_16466_),
    .X(_16666_));
 sky130_fd_sc_hd__nand3_4 _39245_ (.A(_16651_),
    .B(_16652_),
    .C(_16658_),
    .Y(_16667_));
 sky130_fd_sc_hd__nand3_4 _39246_ (.A(_16665_),
    .B(_16666_),
    .C(_16667_),
    .Y(_16668_));
 sky130_fd_sc_hd__and4_1 _39247_ (.A(_19849_),
    .B(_19852_),
    .C(_13456_),
    .D(_13451_),
    .X(_16669_));
 sky130_vsdinv _39248_ (.A(_19848_),
    .Y(_16670_));
 sky130_fd_sc_hd__o22a_1 _39249_ (.A1(_16670_),
    .A2(_11557_),
    .B1(_15009_),
    .B2(_10781_),
    .X(_16671_));
 sky130_fd_sc_hd__or4_4 _39250_ (.A(_08615_),
    .B(_12297_),
    .C(_16669_),
    .D(_16671_),
    .X(_16672_));
 sky130_fd_sc_hd__nor2_1 _39251_ (.A(_16669_),
    .B(_16671_),
    .Y(_16673_));
 sky130_fd_sc_hd__a21o_2 _39252_ (.A1(_19856_),
    .A2(_20089_),
    .B1(_16673_),
    .X(_16674_));
 sky130_fd_sc_hd__o21bai_4 _39253_ (.A1(_16457_),
    .A2(_16455_),
    .B1_N(_16460_),
    .Y(_16675_));
 sky130_fd_sc_hd__a21o_2 _39254_ (.A1(_16672_),
    .A2(_16674_),
    .B1(_16675_),
    .X(_16676_));
 sky130_fd_sc_hd__nand3_4 _39255_ (.A(_16672_),
    .B(_16674_),
    .C(_16675_),
    .Y(_16677_));
 sky130_fd_sc_hd__nand2_4 _39256_ (.A(_16478_),
    .B(_16479_),
    .Y(_16678_));
 sky130_fd_sc_hd__and3_1 _39257_ (.A(_16676_),
    .B(_16677_),
    .C(_16678_),
    .X(_16679_));
 sky130_fd_sc_hd__a21oi_2 _39258_ (.A1(_16676_),
    .A2(_16677_),
    .B1(_16678_),
    .Y(_16680_));
 sky130_fd_sc_hd__o2bb2ai_4 _39259_ (.A1_N(_16664_),
    .A2_N(_16668_),
    .B1(_16679_),
    .B2(_16680_),
    .Y(_16681_));
 sky130_fd_sc_hd__a21oi_4 _39260_ (.A1(_16672_),
    .A2(_16674_),
    .B1(_16675_),
    .Y(_16682_));
 sky130_fd_sc_hd__and3_1 _39261_ (.A(_16672_),
    .B(_16674_),
    .C(_16675_),
    .X(_16683_));
 sky130_fd_sc_hd__o21ai_2 _39262_ (.A1(_16682_),
    .A2(_16683_),
    .B1(_16678_),
    .Y(_16684_));
 sky130_vsdinv _39263_ (.A(_16678_),
    .Y(_16685_));
 sky130_fd_sc_hd__nand3_4 _39264_ (.A(_16676_),
    .B(_16677_),
    .C(_16685_),
    .Y(_16686_));
 sky130_fd_sc_hd__nand2_1 _39265_ (.A(_16684_),
    .B(_16686_),
    .Y(_16687_));
 sky130_fd_sc_hd__nand3_4 _39266_ (.A(_16687_),
    .B(_16668_),
    .C(_16664_),
    .Y(_16688_));
 sky130_fd_sc_hd__nand2_1 _39267_ (.A(_16489_),
    .B(_16488_),
    .Y(_16689_));
 sky130_fd_sc_hd__nand2_4 _39268_ (.A(_16689_),
    .B(_16472_),
    .Y(_16690_));
 sky130_fd_sc_hd__a21oi_4 _39269_ (.A1(_16681_),
    .A2(_16688_),
    .B1(_16690_),
    .Y(_16691_));
 sky130_fd_sc_hd__and3_1 _39270_ (.A(_16681_),
    .B(_16690_),
    .C(_16688_),
    .X(_16692_));
 sky130_fd_sc_hd__nand2_4 _39271_ (.A(_10433_),
    .B(_10259_),
    .Y(_16693_));
 sky130_fd_sc_hd__nand2_4 _39272_ (.A(_07965_),
    .B(_10256_),
    .Y(_16694_));
 sky130_fd_sc_hd__nor2_2 _39273_ (.A(_16693_),
    .B(_16694_),
    .Y(_16695_));
 sky130_fd_sc_hd__nand2_2 _39274_ (.A(_19867_),
    .B(_20074_),
    .Y(_16696_));
 sky130_fd_sc_hd__and2_1 _39275_ (.A(_16693_),
    .B(_16694_),
    .X(_16697_));
 sky130_fd_sc_hd__or3_4 _39276_ (.A(_16695_),
    .B(_16696_),
    .C(_16697_),
    .X(_16698_));
 sky130_fd_sc_hd__o21ai_4 _39277_ (.A1(_16695_),
    .A2(_16697_),
    .B1(_16696_),
    .Y(_16699_));
 sky130_fd_sc_hd__o21bai_4 _39278_ (.A1(_16498_),
    .A2(_16502_),
    .B1_N(_16501_),
    .Y(_16700_));
 sky130_fd_sc_hd__a21oi_4 _39279_ (.A1(_16698_),
    .A2(_16699_),
    .B1(_16700_),
    .Y(_16701_));
 sky130_fd_sc_hd__and3_1 _39280_ (.A(_16698_),
    .B(_16700_),
    .C(_16699_),
    .X(_16702_));
 sky130_fd_sc_hd__and4_1 _39281_ (.A(_18687_),
    .B(_19871_),
    .C(_19875_),
    .D(_20070_),
    .X(_16703_));
 sky130_fd_sc_hd__nand2_2 _39282_ (.A(_14806_),
    .B(_07973_),
    .Y(_16704_));
 sky130_fd_sc_hd__o21a_1 _39283_ (.A1(_16512_),
    .A2(_16147_),
    .B1(_16704_),
    .X(_16705_));
 sky130_fd_sc_hd__nor2_1 _39284_ (.A(_16703_),
    .B(_16705_),
    .Y(_16706_));
 sky130_fd_sc_hd__nor2_1 _39285_ (.A(_16510_),
    .B(_16706_),
    .Y(_16707_));
 sky130_fd_sc_hd__and2_1 _39286_ (.A(_16706_),
    .B(_16510_),
    .X(_16708_));
 sky130_fd_sc_hd__or2_1 _39287_ (.A(_16707_),
    .B(_16708_),
    .X(_16709_));
 sky130_fd_sc_hd__o21ai_4 _39288_ (.A1(_16701_),
    .A2(_16702_),
    .B1(_16709_),
    .Y(_16710_));
 sky130_fd_sc_hd__nor2_2 _39289_ (.A(_16707_),
    .B(_16708_),
    .Y(_16711_));
 sky130_fd_sc_hd__nand3_4 _39290_ (.A(_16698_),
    .B(_16700_),
    .C(_16699_),
    .Y(_16712_));
 sky130_fd_sc_hd__nand3b_4 _39291_ (.A_N(_16701_),
    .B(_16711_),
    .C(_16712_),
    .Y(_16713_));
 sky130_fd_sc_hd__a21oi_2 _39292_ (.A1(_16478_),
    .A2(_16480_),
    .B1(_16481_),
    .Y(_16714_));
 sky130_fd_sc_hd__o21ai_4 _39293_ (.A1(_16485_),
    .A2(_16714_),
    .B1(_16483_),
    .Y(_16715_));
 sky130_fd_sc_hd__a21o_1 _39294_ (.A1(_16710_),
    .A2(_16713_),
    .B1(_16715_),
    .X(_16716_));
 sky130_fd_sc_hd__nand3_4 _39295_ (.A(_16710_),
    .B(_16715_),
    .C(_16713_),
    .Y(_16717_));
 sky130_fd_sc_hd__nand2_2 _39296_ (.A(_16521_),
    .B(_16507_),
    .Y(_16718_));
 sky130_fd_sc_hd__and2_1 _39297_ (.A(_16717_),
    .B(_16718_),
    .X(_16719_));
 sky130_fd_sc_hd__a21oi_4 _39298_ (.A1(_16716_),
    .A2(_16717_),
    .B1(_16718_),
    .Y(_16720_));
 sky130_fd_sc_hd__a21o_2 _39299_ (.A1(_16716_),
    .A2(_16719_),
    .B1(_16720_),
    .X(_16721_));
 sky130_fd_sc_hd__o21ai_4 _39300_ (.A1(_16691_),
    .A2(_16692_),
    .B1(_16721_),
    .Y(_16722_));
 sky130_vsdinv _39301_ (.A(_16489_),
    .Y(_16723_));
 sky130_fd_sc_hd__o21a_1 _39302_ (.A1(_16486_),
    .A2(_16487_),
    .B1(_16472_),
    .X(_16724_));
 sky130_fd_sc_hd__o2bb2ai_4 _39303_ (.A1_N(_16688_),
    .A2_N(_16681_),
    .B1(_16723_),
    .B2(_16724_),
    .Y(_16725_));
 sky130_fd_sc_hd__nand3_1 _39304_ (.A(_16716_),
    .B(_16717_),
    .C(_16718_),
    .Y(_16726_));
 sky130_vsdinv _39305_ (.A(_16726_),
    .Y(_16727_));
 sky130_fd_sc_hd__nor2_4 _39306_ (.A(_16720_),
    .B(_16727_),
    .Y(_16728_));
 sky130_fd_sc_hd__nand3_4 _39307_ (.A(_16681_),
    .B(_16690_),
    .C(_16688_),
    .Y(_16729_));
 sky130_fd_sc_hd__nand3_4 _39308_ (.A(_16725_),
    .B(_16728_),
    .C(_16729_),
    .Y(_16730_));
 sky130_vsdinv _39309_ (.A(_16490_),
    .Y(_16731_));
 sky130_fd_sc_hd__o21ai_2 _39310_ (.A1(_16443_),
    .A2(_16445_),
    .B1(_16491_),
    .Y(_16732_));
 sky130_fd_sc_hd__o2bb2ai_4 _39311_ (.A1_N(_16497_),
    .A2_N(_16532_),
    .B1(_16731_),
    .B2(_16732_),
    .Y(_16733_));
 sky130_fd_sc_hd__a21oi_4 _39312_ (.A1(_16722_),
    .A2(_16730_),
    .B1(_16733_),
    .Y(_16734_));
 sky130_fd_sc_hd__nand2_2 _39313_ (.A(_16497_),
    .B(_16532_),
    .Y(_16735_));
 sky130_fd_sc_hd__nor2_2 _39314_ (.A(_16721_),
    .B(_16691_),
    .Y(_16736_));
 sky130_fd_sc_hd__a21oi_4 _39315_ (.A1(_16725_),
    .A2(_16729_),
    .B1(_16728_),
    .Y(_16737_));
 sky130_fd_sc_hd__a221oi_2 _39316_ (.A1(_16735_),
    .A2(_16492_),
    .B1(_16736_),
    .B2(_16729_),
    .C1(_16737_),
    .Y(_16738_));
 sky130_fd_sc_hd__nand2_1 _39317_ (.A(_16524_),
    .B(_16528_),
    .Y(_16739_));
 sky130_fd_sc_hd__nand2_4 _39318_ (.A(_16739_),
    .B(_16526_),
    .Y(_16740_));
 sky130_fd_sc_hd__o21a_1 _39319_ (.A1(_16549_),
    .A2(_16547_),
    .B1(_16543_),
    .X(_16741_));
 sky130_fd_sc_hd__a21o_1 _39320_ (.A1(_16515_),
    .A2(_16510_),
    .B1(_16511_),
    .X(_16742_));
 sky130_fd_sc_hd__a21o_1 _39321_ (.A1(_16366_),
    .A2(_16364_),
    .B1(_16742_),
    .X(_16743_));
 sky130_fd_sc_hd__nand2_4 _39322_ (.A(_16368_),
    .B(_16742_),
    .Y(_16744_));
 sky130_fd_sc_hd__a21o_1 _39323_ (.A1(_16743_),
    .A2(_16744_),
    .B1(_16545_),
    .X(_16745_));
 sky130_fd_sc_hd__nand3_4 _39324_ (.A(_16743_),
    .B(_16744_),
    .C(_16545_),
    .Y(_16746_));
 sky130_fd_sc_hd__nand3b_4 _39325_ (.A_N(_16741_),
    .B(_16745_),
    .C(_16746_),
    .Y(_16747_));
 sky130_fd_sc_hd__nand2_1 _39326_ (.A(_16745_),
    .B(_16746_),
    .Y(_16748_));
 sky130_fd_sc_hd__nand2_4 _39327_ (.A(_16748_),
    .B(_16741_),
    .Y(_16749_));
 sky130_fd_sc_hd__nand2_1 _39328_ (.A(_16747_),
    .B(_16749_),
    .Y(_16750_));
 sky130_fd_sc_hd__nand2_1 _39329_ (.A(_16750_),
    .B(_16387_),
    .Y(_16751_));
 sky130_fd_sc_hd__nand3_2 _39330_ (.A(_16747_),
    .B(_16749_),
    .C(_16389_),
    .Y(_16752_));
 sky130_fd_sc_hd__nand3b_4 _39331_ (.A_N(_16740_),
    .B(_16751_),
    .C(_16752_),
    .Y(_16753_));
 sky130_fd_sc_hd__nand2_2 _39332_ (.A(_16750_),
    .B(_16389_),
    .Y(_16754_));
 sky130_fd_sc_hd__nand3_4 _39333_ (.A(_16747_),
    .B(_16749_),
    .C(_16387_),
    .Y(_16755_));
 sky130_fd_sc_hd__and2_1 _39334_ (.A(_16557_),
    .B(_16552_),
    .X(_16756_));
 sky130_fd_sc_hd__a31oi_4 _39335_ (.A1(_16754_),
    .A2(_16755_),
    .A3(_16740_),
    .B1(_16756_),
    .Y(_16757_));
 sky130_fd_sc_hd__nand3_4 _39336_ (.A(_16754_),
    .B(_16755_),
    .C(_16740_),
    .Y(_16758_));
 sky130_fd_sc_hd__nand2_2 _39337_ (.A(_16557_),
    .B(_16552_),
    .Y(_16759_));
 sky130_fd_sc_hd__a21oi_4 _39338_ (.A1(_16753_),
    .A2(_16758_),
    .B1(_16759_),
    .Y(_16760_));
 sky130_fd_sc_hd__a21oi_4 _39339_ (.A1(_16753_),
    .A2(_16757_),
    .B1(_16760_),
    .Y(_16761_));
 sky130_fd_sc_hd__o21ai_2 _39340_ (.A1(_16734_),
    .A2(_16738_),
    .B1(_16761_),
    .Y(_16762_));
 sky130_fd_sc_hd__a21boi_4 _39341_ (.A1(_16539_),
    .A2(_16574_),
    .B1_N(_16534_),
    .Y(_16763_));
 sky130_fd_sc_hd__and3_1 _39342_ (.A(_16725_),
    .B(_16728_),
    .C(_16729_),
    .X(_16764_));
 sky130_fd_sc_hd__o21bai_4 _39343_ (.A1(_16737_),
    .A2(_16764_),
    .B1_N(_16733_),
    .Y(_16765_));
 sky130_fd_sc_hd__nand2_1 _39344_ (.A(_16753_),
    .B(_16758_),
    .Y(_16766_));
 sky130_fd_sc_hd__nand2_1 _39345_ (.A(_16766_),
    .B(_16756_),
    .Y(_16767_));
 sky130_fd_sc_hd__nand3_4 _39346_ (.A(_16753_),
    .B(_16758_),
    .C(_16759_),
    .Y(_16768_));
 sky130_fd_sc_hd__nand2_2 _39347_ (.A(_16767_),
    .B(_16768_),
    .Y(_16769_));
 sky130_fd_sc_hd__nand3_4 _39348_ (.A(_16722_),
    .B(_16733_),
    .C(_16730_),
    .Y(_16770_));
 sky130_fd_sc_hd__nand3_4 _39349_ (.A(_16765_),
    .B(_16769_),
    .C(_16770_),
    .Y(_16771_));
 sky130_fd_sc_hd__nand3_4 _39350_ (.A(_16762_),
    .B(_16763_),
    .C(_16771_),
    .Y(_16772_));
 sky130_vsdinv _39351_ (.A(_16768_),
    .Y(_16773_));
 sky130_fd_sc_hd__o22ai_4 _39352_ (.A1(_16760_),
    .A2(_16773_),
    .B1(_16734_),
    .B2(_16738_),
    .Y(_16774_));
 sky130_fd_sc_hd__nand3_4 _39353_ (.A(_16765_),
    .B(_16761_),
    .C(_16770_),
    .Y(_16775_));
 sky130_fd_sc_hd__nand2_1 _39354_ (.A(_16560_),
    .B(_16564_),
    .Y(_16776_));
 sky130_fd_sc_hd__nand2_1 _39355_ (.A(_16776_),
    .B(_16571_),
    .Y(_16777_));
 sky130_fd_sc_hd__nand2_1 _39356_ (.A(_16777_),
    .B(_16568_),
    .Y(_16778_));
 sky130_fd_sc_hd__a21oi_2 _39357_ (.A1(_16531_),
    .A2(_16533_),
    .B1(_16442_),
    .Y(_16779_));
 sky130_fd_sc_hd__o21ai_2 _39358_ (.A1(_16778_),
    .A2(_16779_),
    .B1(_16534_),
    .Y(_16780_));
 sky130_fd_sc_hd__nand3_4 _39359_ (.A(_16774_),
    .B(_16775_),
    .C(_16780_),
    .Y(_16781_));
 sky130_fd_sc_hd__a21o_4 _39360_ (.A1(_16568_),
    .A2(_16560_),
    .B1(_16258_),
    .X(_16782_));
 sky130_fd_sc_hd__buf_4 _39361_ (.A(_16256_),
    .X(_16783_));
 sky130_fd_sc_hd__nor2_4 _39362_ (.A(_16783_),
    .B(_16572_),
    .Y(_16784_));
 sky130_fd_sc_hd__a21oi_4 _39363_ (.A1(_16784_),
    .A2(_16568_),
    .B1(_16587_),
    .Y(_16785_));
 sky130_fd_sc_hd__nand2_2 _39364_ (.A(_16784_),
    .B(_16568_),
    .Y(_16786_));
 sky130_fd_sc_hd__buf_4 _39365_ (.A(_16588_),
    .X(_16787_));
 sky130_fd_sc_hd__a21oi_4 _39366_ (.A1(_16782_),
    .A2(_16786_),
    .B1(_16787_),
    .Y(_16788_));
 sky130_fd_sc_hd__a21oi_4 _39367_ (.A1(_16782_),
    .A2(_16785_),
    .B1(_16788_),
    .Y(_16789_));
 sky130_fd_sc_hd__nand3_4 _39368_ (.A(_16772_),
    .B(_16781_),
    .C(_16789_),
    .Y(_16790_));
 sky130_fd_sc_hd__nand2_2 _39369_ (.A(_16785_),
    .B(_16782_),
    .Y(_16791_));
 sky130_vsdinv _39370_ (.A(_16791_),
    .Y(_16792_));
 sky130_fd_sc_hd__o2bb2ai_4 _39371_ (.A1_N(_16781_),
    .A2_N(_16772_),
    .B1(_16788_),
    .B2(_16792_),
    .Y(_16793_));
 sky130_fd_sc_hd__o211a_4 _39372_ (.A1(_16584_),
    .A2(_16643_),
    .B1(_16790_),
    .C1(_16793_),
    .X(_16794_));
 sky130_fd_sc_hd__nand2_1 _39373_ (.A(_16793_),
    .B(_16790_),
    .Y(_16795_));
 sky130_fd_sc_hd__nor2_1 _39374_ (.A(_16584_),
    .B(_16643_),
    .Y(_16796_));
 sky130_fd_sc_hd__nand2_2 _39375_ (.A(_16795_),
    .B(_16796_),
    .Y(_16797_));
 sky130_fd_sc_hd__nand2_2 _39376_ (.A(_16589_),
    .B(_16590_),
    .Y(_16798_));
 sky130_fd_sc_hd__nor2_8 _39377_ (.A(_14354_),
    .B(_16798_),
    .Y(_16799_));
 sky130_vsdinv _39378_ (.A(_16798_),
    .Y(_16800_));
 sky130_fd_sc_hd__nor2_8 _39379_ (.A(_14931_),
    .B(_16800_),
    .Y(_16801_));
 sky130_fd_sc_hd__nor2_8 _39380_ (.A(_16799_),
    .B(_16801_),
    .Y(_16802_));
 sky130_vsdinv _39381_ (.A(_16802_),
    .Y(_16803_));
 sky130_fd_sc_hd__nand2_1 _39382_ (.A(_16797_),
    .B(_16803_),
    .Y(_16804_));
 sky130_fd_sc_hd__o21ai_4 _39383_ (.A1(_16594_),
    .A2(_16578_),
    .B1(_16602_),
    .Y(_16805_));
 sky130_fd_sc_hd__a21oi_4 _39384_ (.A1(_16793_),
    .A2(_16790_),
    .B1(_16805_),
    .Y(_16806_));
 sky130_fd_sc_hd__o21ai_2 _39385_ (.A1(_16806_),
    .A2(_16794_),
    .B1(_16802_),
    .Y(_16807_));
 sky130_fd_sc_hd__nand2_1 _39386_ (.A(_16409_),
    .B(_16411_),
    .Y(_16808_));
 sky130_fd_sc_hd__a22oi_4 _39387_ (.A1(_16410_),
    .A2(_16808_),
    .B1(_16605_),
    .B2(_16607_),
    .Y(_16809_));
 sky130_fd_sc_hd__a21o_1 _39388_ (.A1(_16608_),
    .A2(_16615_),
    .B1(_16809_),
    .X(_16810_));
 sky130_fd_sc_hd__o211ai_4 _39389_ (.A1(_16794_),
    .A2(_16804_),
    .B1(_16807_),
    .C1(_16810_),
    .Y(_16811_));
 sky130_fd_sc_hd__o22ai_4 _39390_ (.A1(_16801_),
    .A2(_16799_),
    .B1(_16806_),
    .B2(_16794_),
    .Y(_16812_));
 sky130_fd_sc_hd__a21oi_2 _39391_ (.A1(_16608_),
    .A2(_16615_),
    .B1(_16809_),
    .Y(_16813_));
 sky130_vsdinv _39392_ (.A(_16790_),
    .Y(_16814_));
 sky130_fd_sc_hd__nand2_2 _39393_ (.A(_16805_),
    .B(_16793_),
    .Y(_16815_));
 sky130_fd_sc_hd__o211ai_4 _39394_ (.A1(_16814_),
    .A2(_16815_),
    .B1(_16802_),
    .C1(_16797_),
    .Y(_16816_));
 sky130_fd_sc_hd__nand3_4 _39395_ (.A(_16812_),
    .B(_16813_),
    .C(_16816_),
    .Y(_16817_));
 sky130_fd_sc_hd__buf_6 _39396_ (.A(net411),
    .X(_16818_));
 sky130_fd_sc_hd__nor2_4 _39397_ (.A(_16818_),
    .B(_16612_),
    .Y(_16819_));
 sky130_fd_sc_hd__a21oi_4 _39398_ (.A1(_16811_),
    .A2(_16817_),
    .B1(_16819_),
    .Y(_16820_));
 sky130_fd_sc_hd__a31oi_4 _39399_ (.A1(_16614_),
    .A2(_16618_),
    .A3(_16616_),
    .B1(_16424_),
    .Y(_16821_));
 sky130_fd_sc_hd__nand3_2 _39400_ (.A(_16811_),
    .B(_16819_),
    .C(_16817_),
    .Y(_16822_));
 sky130_fd_sc_hd__o21ai_4 _39401_ (.A1(_16619_),
    .A2(_16821_),
    .B1(_16822_),
    .Y(_16823_));
 sky130_vsdinv _39402_ (.A(_16819_),
    .Y(_16824_));
 sky130_fd_sc_hd__a21o_1 _39403_ (.A1(_16811_),
    .A2(_16817_),
    .B1(_16824_),
    .X(_16825_));
 sky130_fd_sc_hd__nand3b_2 _39404_ (.A_N(_16819_),
    .B(_16811_),
    .C(_16817_),
    .Y(_16826_));
 sky130_fd_sc_hd__nor2_2 _39405_ (.A(_16619_),
    .B(_16821_),
    .Y(_16827_));
 sky130_fd_sc_hd__nand3_4 _39406_ (.A(_16825_),
    .B(_16826_),
    .C(_16827_),
    .Y(_16828_));
 sky130_fd_sc_hd__o21a_1 _39407_ (.A1(_16820_),
    .A2(_16823_),
    .B1(_16828_),
    .X(_16829_));
 sky130_vsdinv _39408_ (.A(_16635_),
    .Y(_16830_));
 sky130_fd_sc_hd__o21ai_1 _39409_ (.A1(_16830_),
    .A2(_16642_),
    .B1(_16631_),
    .Y(_16831_));
 sky130_fd_sc_hd__xor2_1 _39410_ (.A(_16829_),
    .B(_16831_),
    .X(_02670_));
 sky130_fd_sc_hd__a21oi_4 _39411_ (.A1(_16797_),
    .A2(_16803_),
    .B1(_16794_),
    .Y(_16832_));
 sky130_fd_sc_hd__nand2_4 _39412_ (.A(_16791_),
    .B(_16782_),
    .Y(_16833_));
 sky130_vsdinv _39413_ (.A(_16833_),
    .Y(_16834_));
 sky130_fd_sc_hd__nor2_8 _39414_ (.A(_16423_),
    .B(_16834_),
    .Y(_16835_));
 sky130_fd_sc_hd__nor2_8 _39415_ (.A(net413),
    .B(_16833_),
    .Y(_16836_));
 sky130_fd_sc_hd__a21oi_1 _39416_ (.A1(_16366_),
    .A2(_16364_),
    .B1(_16742_),
    .Y(_16837_));
 sky130_fd_sc_hd__o21ai_2 _39417_ (.A1(_16549_),
    .A2(_16837_),
    .B1(_16744_),
    .Y(_16838_));
 sky130_fd_sc_hd__o21bai_4 _39418_ (.A1(_16509_),
    .A2(_16705_),
    .B1_N(_16703_),
    .Y(_16839_));
 sky130_fd_sc_hd__nand2_1 _39419_ (.A(_16365_),
    .B(_15813_),
    .Y(_16840_));
 sky130_fd_sc_hd__nand2_4 _39420_ (.A(_16361_),
    .B(net456),
    .Y(_16841_));
 sky130_fd_sc_hd__and2_2 _39421_ (.A(_16840_),
    .B(_16841_),
    .X(_16842_));
 sky130_fd_sc_hd__xor2_4 _39422_ (.A(_16839_),
    .B(_16842_),
    .X(_16843_));
 sky130_fd_sc_hd__nand2_4 _39423_ (.A(_16838_),
    .B(_16843_),
    .Y(_16844_));
 sky130_fd_sc_hd__xnor2_2 _39424_ (.A(_16839_),
    .B(_16842_),
    .Y(_16845_));
 sky130_fd_sc_hd__nand3_4 _39425_ (.A(_16746_),
    .B(_16744_),
    .C(_16845_),
    .Y(_16846_));
 sky130_fd_sc_hd__a21oi_2 _39426_ (.A1(_16844_),
    .A2(_16846_),
    .B1(_16170_),
    .Y(_16847_));
 sky130_fd_sc_hd__and3_1 _39427_ (.A(_16844_),
    .B(_16846_),
    .C(_15840_),
    .X(_16848_));
 sky130_fd_sc_hd__a21oi_4 _39428_ (.A1(_16710_),
    .A2(_16713_),
    .B1(_16715_),
    .Y(_16849_));
 sky130_vsdinv _39429_ (.A(_16718_),
    .Y(_16850_));
 sky130_fd_sc_hd__o21ai_4 _39430_ (.A1(_16849_),
    .A2(_16850_),
    .B1(_16717_),
    .Y(_16851_));
 sky130_fd_sc_hd__o21ai_4 _39431_ (.A1(_16847_),
    .A2(_16848_),
    .B1(_16851_),
    .Y(_16852_));
 sky130_fd_sc_hd__nand3_4 _39432_ (.A(_16844_),
    .B(_16846_),
    .C(_16170_),
    .Y(_16853_));
 sky130_fd_sc_hd__a21o_1 _39433_ (.A1(_16844_),
    .A2(_16846_),
    .B1(_15840_),
    .X(_16854_));
 sky130_fd_sc_hd__o2111ai_4 _39434_ (.A1(_16849_),
    .A2(_16850_),
    .B1(_16717_),
    .C1(_16853_),
    .D1(_16854_),
    .Y(_16855_));
 sky130_fd_sc_hd__nand2_2 _39435_ (.A(_16749_),
    .B(_16172_),
    .Y(_16856_));
 sky130_fd_sc_hd__nand2_2 _39436_ (.A(_16856_),
    .B(_16747_),
    .Y(_16857_));
 sky130_fd_sc_hd__a21oi_4 _39437_ (.A1(_16852_),
    .A2(_16855_),
    .B1(_16857_),
    .Y(_16858_));
 sky130_fd_sc_hd__and3_1 _39438_ (.A(_16852_),
    .B(_16857_),
    .C(_16855_),
    .X(_16859_));
 sky130_fd_sc_hd__nand2_4 _39439_ (.A(_19868_),
    .B(_10779_),
    .Y(_16860_));
 sky130_fd_sc_hd__nand2_2 _39440_ (.A(_10440_),
    .B(_11587_),
    .Y(_16861_));
 sky130_fd_sc_hd__nand2_4 _39441_ (.A(_08592_),
    .B(_11173_),
    .Y(_16862_));
 sky130_fd_sc_hd__nor2_1 _39442_ (.A(_16861_),
    .B(_16862_),
    .Y(_16863_));
 sky130_fd_sc_hd__and2_1 _39443_ (.A(_16861_),
    .B(_16862_),
    .X(_16864_));
 sky130_fd_sc_hd__or2_2 _39444_ (.A(_16863_),
    .B(_16864_),
    .X(_16865_));
 sky130_fd_sc_hd__or2_4 _39445_ (.A(_16860_),
    .B(_16865_),
    .X(_16866_));
 sky130_fd_sc_hd__nand2_4 _39446_ (.A(_16865_),
    .B(_16860_),
    .Y(_16867_));
 sky130_fd_sc_hd__o21ai_4 _39447_ (.A1(_16693_),
    .A2(_16694_),
    .B1(_16698_),
    .Y(_16868_));
 sky130_fd_sc_hd__a21oi_4 _39448_ (.A1(_16866_),
    .A2(_16867_),
    .B1(_16868_),
    .Y(_16869_));
 sky130_fd_sc_hd__nor2_1 _39449_ (.A(_16860_),
    .B(_16865_),
    .Y(_16870_));
 sky130_fd_sc_hd__and3b_2 _39450_ (.A_N(_16870_),
    .B(_16868_),
    .C(_16867_),
    .X(_16871_));
 sky130_fd_sc_hd__nand2_2 _39451_ (.A(_14806_),
    .B(_10628_),
    .Y(_16872_));
 sky130_fd_sc_hd__or2_1 _39452_ (.A(_16704_),
    .B(_16872_),
    .X(_16873_));
 sky130_fd_sc_hd__nand2_1 _39453_ (.A(_16704_),
    .B(_16872_),
    .Y(_16874_));
 sky130_fd_sc_hd__nand2_1 _39454_ (.A(_16873_),
    .B(_16874_),
    .Y(_16875_));
 sky130_fd_sc_hd__or2_2 _39455_ (.A(_16509_),
    .B(_16875_),
    .X(_16876_));
 sky130_fd_sc_hd__nand2_1 _39456_ (.A(_16875_),
    .B(_16509_),
    .Y(_16877_));
 sky130_fd_sc_hd__and2_2 _39457_ (.A(_16876_),
    .B(_16877_),
    .X(_16878_));
 sky130_fd_sc_hd__clkbuf_4 _39458_ (.A(_16878_),
    .X(_16879_));
 sky130_fd_sc_hd__o21ai_2 _39459_ (.A1(_16869_),
    .A2(_16871_),
    .B1(_16879_),
    .Y(_16880_));
 sky130_fd_sc_hd__a21oi_4 _39460_ (.A1(_16676_),
    .A2(_16678_),
    .B1(_16683_),
    .Y(_16881_));
 sky130_fd_sc_hd__a21o_2 _39461_ (.A1(_16866_),
    .A2(_16867_),
    .B1(_16868_),
    .X(_16882_));
 sky130_fd_sc_hd__nand3_4 _39462_ (.A(_16866_),
    .B(_16868_),
    .C(_16867_),
    .Y(_16883_));
 sky130_fd_sc_hd__nand2_4 _39463_ (.A(_16876_),
    .B(_16877_),
    .Y(_16884_));
 sky130_fd_sc_hd__buf_4 _39464_ (.A(_16884_),
    .X(_16885_));
 sky130_fd_sc_hd__nand3_2 _39465_ (.A(_16882_),
    .B(_16883_),
    .C(_16885_),
    .Y(_16886_));
 sky130_fd_sc_hd__nand3_4 _39466_ (.A(_16880_),
    .B(_16881_),
    .C(_16886_),
    .Y(_16887_));
 sky130_fd_sc_hd__o21ai_2 _39467_ (.A1(_16869_),
    .A2(_16871_),
    .B1(_16884_),
    .Y(_16888_));
 sky130_fd_sc_hd__o21ai_4 _39468_ (.A1(_16685_),
    .A2(_16682_),
    .B1(_16677_),
    .Y(_16889_));
 sky130_fd_sc_hd__nand3_4 _39469_ (.A(_16882_),
    .B(_16883_),
    .C(_16878_),
    .Y(_16890_));
 sky130_fd_sc_hd__nand3_4 _39470_ (.A(_16888_),
    .B(_16889_),
    .C(_16890_),
    .Y(_16891_));
 sky130_fd_sc_hd__nand2_4 _39471_ (.A(_16713_),
    .B(_16712_),
    .Y(_16892_));
 sky130_fd_sc_hd__a21oi_4 _39472_ (.A1(_16887_),
    .A2(_16891_),
    .B1(_16892_),
    .Y(_16893_));
 sky130_fd_sc_hd__nand3_4 _39473_ (.A(_16887_),
    .B(_16891_),
    .C(_16892_),
    .Y(_16894_));
 sky130_vsdinv _39474_ (.A(_16894_),
    .Y(_16895_));
 sky130_fd_sc_hd__nor2_4 _39475_ (.A(_10405_),
    .B(_12100_),
    .Y(_16896_));
 sky130_fd_sc_hd__and4_2 _39476_ (.A(_10824_),
    .B(_18695_),
    .C(_15907_),
    .D(_13758_),
    .X(_16897_));
 sky130_fd_sc_hd__o22a_2 _39477_ (.A1(_20112_),
    .A2(_15914_),
    .B1(_16103_),
    .B2(_12093_),
    .X(_16898_));
 sky130_fd_sc_hd__or3_4 _39478_ (.A(_16896_),
    .B(_16897_),
    .C(_16898_),
    .X(_16899_));
 sky130_fd_sc_hd__o21ai_4 _39479_ (.A1(_16897_),
    .A2(_16898_),
    .B1(_16896_),
    .Y(_16900_));
 sky130_fd_sc_hd__nor2_1 _39480_ (.A(_16644_),
    .B(_16645_),
    .Y(_16901_));
 sky130_fd_sc_hd__or2_4 _39481_ (.A(_16646_),
    .B(_16901_),
    .X(_16902_));
 sky130_fd_sc_hd__a21o_1 _39482_ (.A1(_16899_),
    .A2(_16900_),
    .B1(_16902_),
    .X(_16903_));
 sky130_fd_sc_hd__nand3_4 _39483_ (.A(_16902_),
    .B(_16900_),
    .C(_16899_),
    .Y(_16904_));
 sky130_fd_sc_hd__nor2_4 _39484_ (.A(_09321_),
    .B(_11563_),
    .Y(_16905_));
 sky130_fd_sc_hd__a22o_1 _39485_ (.A1(_19837_),
    .A2(_20103_),
    .B1(_19842_),
    .B2(_20099_),
    .X(_16906_));
 sky130_fd_sc_hd__o21ai_4 _39486_ (.A1(_16311_),
    .A2(_11737_),
    .B1(_16906_),
    .Y(_16907_));
 sky130_fd_sc_hd__xnor2_4 _39487_ (.A(_16905_),
    .B(_16907_),
    .Y(_16908_));
 sky130_fd_sc_hd__a21o_1 _39488_ (.A1(_16903_),
    .A2(_16904_),
    .B1(_16908_),
    .X(_16909_));
 sky130_fd_sc_hd__a21oi_2 _39489_ (.A1(_16647_),
    .A2(_16648_),
    .B1(_16650_),
    .Y(_16910_));
 sky130_fd_sc_hd__a21o_1 _39490_ (.A1(_16662_),
    .A2(_16652_),
    .B1(_16910_),
    .X(_16911_));
 sky130_fd_sc_hd__nand3_2 _39491_ (.A(_16903_),
    .B(_16904_),
    .C(_16908_),
    .Y(_16912_));
 sky130_fd_sc_hd__nand3_4 _39492_ (.A(_16909_),
    .B(_16911_),
    .C(_16912_),
    .Y(_16913_));
 sky130_fd_sc_hd__a21oi_4 _39493_ (.A1(_16899_),
    .A2(_16900_),
    .B1(_16902_),
    .Y(_16914_));
 sky130_fd_sc_hd__and3_1 _39494_ (.A(_16902_),
    .B(_16899_),
    .C(_16900_),
    .X(_16915_));
 sky130_fd_sc_hd__o21ai_2 _39495_ (.A1(_16914_),
    .A2(_16915_),
    .B1(_16908_),
    .Y(_16916_));
 sky130_fd_sc_hd__a21oi_2 _39496_ (.A1(_16662_),
    .A2(_16652_),
    .B1(_16910_),
    .Y(_16917_));
 sky130_fd_sc_hd__nand3b_2 _39497_ (.A_N(_16908_),
    .B(_16903_),
    .C(_16904_),
    .Y(_16918_));
 sky130_fd_sc_hd__nand3_4 _39498_ (.A(_16916_),
    .B(_16917_),
    .C(_16918_),
    .Y(_16919_));
 sky130_fd_sc_hd__nand2_1 _39499_ (.A(_19849_),
    .B(_13456_),
    .Y(_16920_));
 sky130_fd_sc_hd__o21a_1 _39500_ (.A1(_15010_),
    .A2(_12297_),
    .B1(_16920_),
    .X(_16921_));
 sky130_fd_sc_hd__or2_1 _39501_ (.A(_16920_),
    .B(_15010_),
    .X(_16922_));
 sky130_fd_sc_hd__nor2_4 _39502_ (.A(_12297_),
    .B(_16922_),
    .Y(_16923_));
 sky130_fd_sc_hd__nand2_1 _39503_ (.A(_19856_),
    .B(_20084_),
    .Y(_16924_));
 sky130_fd_sc_hd__o21ai_1 _39504_ (.A1(_16921_),
    .A2(_16923_),
    .B1(_16924_),
    .Y(_16925_));
 sky130_fd_sc_hd__nor2_1 _39505_ (.A(_16920_),
    .B(_15010_),
    .Y(_16926_));
 sky130_fd_sc_hd__a211o_1 _39506_ (.A1(_20089_),
    .A2(_16926_),
    .B1(_16924_),
    .C1(_16921_),
    .X(_16927_));
 sky130_fd_sc_hd__a32o_1 _39507_ (.A1(_16093_),
    .A2(_20103_),
    .A3(_20106_),
    .B1(_16656_),
    .B2(_16655_),
    .X(_16928_));
 sky130_fd_sc_hd__a21o_1 _39508_ (.A1(_16925_),
    .A2(_16927_),
    .B1(_16928_),
    .X(_16929_));
 sky130_fd_sc_hd__nand3_2 _39509_ (.A(_16925_),
    .B(_16928_),
    .C(_16927_),
    .Y(_16930_));
 sky130_fd_sc_hd__a31o_1 _39510_ (.A1(_16673_),
    .A2(_19856_),
    .A3(_20089_),
    .B1(_16669_),
    .X(_16931_));
 sky130_vsdinv _39511_ (.A(_16931_),
    .Y(_16932_));
 sky130_fd_sc_hd__a21o_1 _39512_ (.A1(_16929_),
    .A2(_16930_),
    .B1(_16932_),
    .X(_16933_));
 sky130_fd_sc_hd__nand3b_1 _39513_ (.A_N(_16931_),
    .B(_16929_),
    .C(_16930_),
    .Y(_16934_));
 sky130_fd_sc_hd__nand2_2 _39514_ (.A(_16933_),
    .B(_16934_),
    .Y(_16935_));
 sky130_fd_sc_hd__a21o_2 _39515_ (.A1(_16913_),
    .A2(_16919_),
    .B1(_16935_),
    .X(_16936_));
 sky130_fd_sc_hd__nand3_4 _39516_ (.A(_16913_),
    .B(_16919_),
    .C(_16935_),
    .Y(_16937_));
 sky130_fd_sc_hd__nand2_2 _39517_ (.A(_16688_),
    .B(_16664_),
    .Y(_16938_));
 sky130_fd_sc_hd__a21oi_4 _39518_ (.A1(_16936_),
    .A2(_16937_),
    .B1(_16938_),
    .Y(_16939_));
 sky130_vsdinv _39519_ (.A(_16664_),
    .Y(_16940_));
 sky130_fd_sc_hd__a32oi_4 _39520_ (.A1(_16665_),
    .A2(_16666_),
    .A3(_16667_),
    .B1(_16686_),
    .B2(_16684_),
    .Y(_16941_));
 sky130_fd_sc_hd__o211a_1 _39521_ (.A1(_16940_),
    .A2(_16941_),
    .B1(_16937_),
    .C1(_16936_),
    .X(_16942_));
 sky130_fd_sc_hd__o22ai_4 _39522_ (.A1(_16893_),
    .A2(_16895_),
    .B1(_16939_),
    .B2(_16942_),
    .Y(_16943_));
 sky130_fd_sc_hd__nand2_1 _39523_ (.A(_16936_),
    .B(_16937_),
    .Y(_16944_));
 sky130_fd_sc_hd__nor2_1 _39524_ (.A(_16940_),
    .B(_16941_),
    .Y(_16945_));
 sky130_fd_sc_hd__nand2_1 _39525_ (.A(_16944_),
    .B(_16945_),
    .Y(_16946_));
 sky130_fd_sc_hd__nand3_4 _39526_ (.A(_16938_),
    .B(_16936_),
    .C(_16937_),
    .Y(_16947_));
 sky130_vsdinv _39527_ (.A(_16892_),
    .Y(_16948_));
 sky130_fd_sc_hd__a31oi_2 _39528_ (.A1(_16888_),
    .A2(_16889_),
    .A3(_16890_),
    .B1(_16948_),
    .Y(_16949_));
 sky130_fd_sc_hd__a21oi_2 _39529_ (.A1(_16949_),
    .A2(_16887_),
    .B1(_16893_),
    .Y(_16950_));
 sky130_fd_sc_hd__nand3_4 _39530_ (.A(_16946_),
    .B(_16947_),
    .C(_16950_),
    .Y(_16951_));
 sky130_fd_sc_hd__o21ai_4 _39531_ (.A1(_16721_),
    .A2(_16691_),
    .B1(_16729_),
    .Y(_16952_));
 sky130_fd_sc_hd__a21oi_4 _39532_ (.A1(_16943_),
    .A2(_16951_),
    .B1(_16952_),
    .Y(_16953_));
 sky130_fd_sc_hd__o211a_2 _39533_ (.A1(_16692_),
    .A2(_16736_),
    .B1(_16951_),
    .C1(_16943_),
    .X(_16954_));
 sky130_fd_sc_hd__o22ai_4 _39534_ (.A1(_16858_),
    .A2(_16859_),
    .B1(_16953_),
    .B2(_16954_),
    .Y(_16955_));
 sky130_fd_sc_hd__o21ai_2 _39535_ (.A1(_16769_),
    .A2(_16734_),
    .B1(_16770_),
    .Y(_16956_));
 sky130_fd_sc_hd__a21o_1 _39536_ (.A1(_16943_),
    .A2(_16951_),
    .B1(_16952_),
    .X(_16957_));
 sky130_fd_sc_hd__nand2_1 _39537_ (.A(_16854_),
    .B(_16853_),
    .Y(_16958_));
 sky130_fd_sc_hd__a22oi_4 _39538_ (.A1(_16856_),
    .A2(_16747_),
    .B1(_16958_),
    .B2(_16851_),
    .Y(_16959_));
 sky130_fd_sc_hd__a21oi_4 _39539_ (.A1(_16855_),
    .A2(_16959_),
    .B1(_16858_),
    .Y(_16960_));
 sky130_fd_sc_hd__nand3_4 _39540_ (.A(_16943_),
    .B(_16952_),
    .C(_16951_),
    .Y(_16961_));
 sky130_fd_sc_hd__nand3_2 _39541_ (.A(_16957_),
    .B(_16960_),
    .C(_16961_),
    .Y(_16962_));
 sky130_fd_sc_hd__nand3_4 _39542_ (.A(_16955_),
    .B(_16956_),
    .C(_16962_),
    .Y(_16963_));
 sky130_fd_sc_hd__o21ai_4 _39543_ (.A1(_16953_),
    .A2(_16954_),
    .B1(_16960_),
    .Y(_16964_));
 sky130_fd_sc_hd__nand2_1 _39544_ (.A(_16725_),
    .B(_16729_),
    .Y(_16965_));
 sky130_fd_sc_hd__a22oi_4 _39545_ (.A1(_16735_),
    .A2(_16492_),
    .B1(_16721_),
    .B2(_16965_),
    .Y(_16966_));
 sky130_fd_sc_hd__a22oi_4 _39546_ (.A1(_16730_),
    .A2(_16966_),
    .B1(_16765_),
    .B2(_16761_),
    .Y(_16967_));
 sky130_fd_sc_hd__a21o_1 _39547_ (.A1(_16855_),
    .A2(_16959_),
    .B1(_16858_),
    .X(_16968_));
 sky130_fd_sc_hd__nand3_4 _39548_ (.A(_16957_),
    .B(_16968_),
    .C(_16961_),
    .Y(_16969_));
 sky130_fd_sc_hd__nand3_4 _39549_ (.A(_16964_),
    .B(_16967_),
    .C(_16969_),
    .Y(_16970_));
 sky130_fd_sc_hd__buf_4 _39550_ (.A(_16257_),
    .X(_16971_));
 sky130_fd_sc_hd__a21o_1 _39551_ (.A1(_16768_),
    .A2(_16758_),
    .B1(_16971_),
    .X(_16972_));
 sky130_fd_sc_hd__nand2_1 _39552_ (.A(_16758_),
    .B(_16257_),
    .Y(_16973_));
 sky130_fd_sc_hd__a21o_1 _39553_ (.A1(_16757_),
    .A2(_16753_),
    .B1(_16973_),
    .X(_16974_));
 sky130_fd_sc_hd__clkbuf_4 _39554_ (.A(_16592_),
    .X(_16975_));
 sky130_fd_sc_hd__a21oi_2 _39555_ (.A1(_16972_),
    .A2(_16974_),
    .B1(_16975_),
    .Y(_16976_));
 sky130_fd_sc_hd__a21oi_4 _39556_ (.A1(_16768_),
    .A2(_16758_),
    .B1(_16971_),
    .Y(_16977_));
 sky130_fd_sc_hd__nand2_2 _39557_ (.A(_16974_),
    .B(_16592_),
    .Y(_16978_));
 sky130_fd_sc_hd__nor2_2 _39558_ (.A(_16977_),
    .B(_16978_),
    .Y(_16979_));
 sky130_fd_sc_hd__o2bb2ai_4 _39559_ (.A1_N(_16963_),
    .A2_N(_16970_),
    .B1(_16976_),
    .B2(_16979_),
    .Y(_16980_));
 sky130_fd_sc_hd__a21oi_1 _39560_ (.A1(_16757_),
    .A2(_16753_),
    .B1(_16973_),
    .Y(_16981_));
 sky130_fd_sc_hd__buf_4 _39561_ (.A(_16587_),
    .X(_16982_));
 sky130_fd_sc_hd__o21ai_1 _39562_ (.A1(_16981_),
    .A2(_16977_),
    .B1(_16982_),
    .Y(_16983_));
 sky130_fd_sc_hd__o21ai_2 _39563_ (.A1(_16977_),
    .A2(_16978_),
    .B1(_16983_),
    .Y(_16984_));
 sky130_vsdinv _39564_ (.A(_16984_),
    .Y(_16985_));
 sky130_fd_sc_hd__nand3_4 _39565_ (.A(_16985_),
    .B(_16970_),
    .C(_16963_),
    .Y(_16986_));
 sky130_fd_sc_hd__nand2_1 _39566_ (.A(_16772_),
    .B(_16789_),
    .Y(_16987_));
 sky130_fd_sc_hd__nand2_4 _39567_ (.A(_16987_),
    .B(_16781_),
    .Y(_16988_));
 sky130_fd_sc_hd__a21oi_4 _39568_ (.A1(_16980_),
    .A2(_16986_),
    .B1(_16988_),
    .Y(_16989_));
 sky130_fd_sc_hd__and3_1 _39569_ (.A(_16774_),
    .B(_16780_),
    .C(_16775_),
    .X(_16990_));
 sky130_fd_sc_hd__nand2_1 _39570_ (.A(_16782_),
    .B(_16786_),
    .Y(_16991_));
 sky130_fd_sc_hd__buf_4 _39571_ (.A(_16587_),
    .X(_16992_));
 sky130_fd_sc_hd__nand2_1 _39572_ (.A(_16991_),
    .B(_16992_),
    .Y(_16993_));
 sky130_fd_sc_hd__nand2_1 _39573_ (.A(_16993_),
    .B(_16791_),
    .Y(_16994_));
 sky130_fd_sc_hd__a31oi_1 _39574_ (.A1(_16762_),
    .A2(_16763_),
    .A3(_16771_),
    .B1(_16994_),
    .Y(_16995_));
 sky130_fd_sc_hd__o211a_2 _39575_ (.A1(_16990_),
    .A2(_16995_),
    .B1(_16986_),
    .C1(_16980_),
    .X(_16996_));
 sky130_fd_sc_hd__o22ai_4 _39576_ (.A1(_16835_),
    .A2(_16836_),
    .B1(_16989_),
    .B2(_16996_),
    .Y(_16997_));
 sky130_fd_sc_hd__a21o_1 _39577_ (.A1(_16980_),
    .A2(_16986_),
    .B1(_16988_),
    .X(_16998_));
 sky130_fd_sc_hd__nand3_4 _39578_ (.A(_16988_),
    .B(_16980_),
    .C(_16986_),
    .Y(_16999_));
 sky130_fd_sc_hd__nor2_8 _39579_ (.A(_16836_),
    .B(_16835_),
    .Y(_17000_));
 sky130_fd_sc_hd__nand3_4 _39580_ (.A(_16998_),
    .B(_16999_),
    .C(_17000_),
    .Y(_17001_));
 sky130_fd_sc_hd__nand3_4 _39581_ (.A(_16832_),
    .B(_16997_),
    .C(_17001_),
    .Y(_17002_));
 sky130_fd_sc_hd__nor2_8 _39582_ (.A(net412),
    .B(_16834_),
    .Y(_17003_));
 sky130_fd_sc_hd__buf_4 _39583_ (.A(_16426_),
    .X(_17004_));
 sky130_fd_sc_hd__nor2_2 _39584_ (.A(_17004_),
    .B(_16833_),
    .Y(_17005_));
 sky130_fd_sc_hd__o22ai_4 _39585_ (.A1(_17003_),
    .A2(_17005_),
    .B1(_16989_),
    .B2(_16996_),
    .Y(_17006_));
 sky130_vsdinv _39586_ (.A(_17000_),
    .Y(_17007_));
 sky130_fd_sc_hd__nand3_4 _39587_ (.A(_16998_),
    .B(_16999_),
    .C(_17007_),
    .Y(_17008_));
 sky130_fd_sc_hd__o22ai_4 _39588_ (.A1(_16814_),
    .A2(_16815_),
    .B1(_16802_),
    .B2(_16806_),
    .Y(_17009_));
 sky130_fd_sc_hd__nand3_4 _39589_ (.A(_17006_),
    .B(_17008_),
    .C(_17009_),
    .Y(_17010_));
 sky130_fd_sc_hd__nor2_4 _39590_ (.A(net411),
    .B(_16800_),
    .Y(_17011_));
 sky130_fd_sc_hd__a21oi_1 _39591_ (.A1(_17002_),
    .A2(_17010_),
    .B1(_17011_),
    .Y(_17012_));
 sky130_fd_sc_hd__and3_1 _39592_ (.A(_17002_),
    .B(_17010_),
    .C(_17011_),
    .X(_17013_));
 sky130_fd_sc_hd__nand2_1 _39593_ (.A(_16817_),
    .B(_16819_),
    .Y(_17014_));
 sky130_fd_sc_hd__nand2_2 _39594_ (.A(_17014_),
    .B(_16811_),
    .Y(_17015_));
 sky130_fd_sc_hd__o21bai_2 _39595_ (.A1(_17012_),
    .A2(_17013_),
    .B1_N(_17015_),
    .Y(_17016_));
 sky130_fd_sc_hd__and3_1 _39596_ (.A(_17006_),
    .B(_17009_),
    .C(_17008_),
    .X(_17017_));
 sky130_fd_sc_hd__nand2_2 _39597_ (.A(_17002_),
    .B(_17011_),
    .Y(_17018_));
 sky130_fd_sc_hd__nand2_1 _39598_ (.A(_17002_),
    .B(_17010_),
    .Y(_17019_));
 sky130_vsdinv _39599_ (.A(_17011_),
    .Y(_17020_));
 sky130_fd_sc_hd__nand2_1 _39600_ (.A(_17019_),
    .B(_17020_),
    .Y(_17021_));
 sky130_fd_sc_hd__o211ai_4 _39601_ (.A1(_17017_),
    .A2(_17018_),
    .B1(_17015_),
    .C1(_17021_),
    .Y(_17022_));
 sky130_fd_sc_hd__and2_1 _39602_ (.A(_17016_),
    .B(_17022_),
    .X(_17023_));
 sky130_fd_sc_hd__o2111a_1 _39603_ (.A1(_16820_),
    .A2(_16823_),
    .B1(_16635_),
    .C1(_16631_),
    .D1(_16828_),
    .X(_17024_));
 sky130_fd_sc_hd__nand2_1 _39604_ (.A(_16632_),
    .B(_16634_),
    .Y(_17025_));
 sky130_fd_sc_hd__nor2_1 _39605_ (.A(_16820_),
    .B(_16823_),
    .Y(_17026_));
 sky130_fd_sc_hd__a31o_1 _39606_ (.A1(_16828_),
    .A2(_17025_),
    .A3(_16624_),
    .B1(_17026_),
    .X(_17027_));
 sky130_fd_sc_hd__a21oi_4 _39607_ (.A1(_17024_),
    .A2(_16641_),
    .B1(_17027_),
    .Y(_17028_));
 sky130_vsdinv _39608_ (.A(_17028_),
    .Y(_17029_));
 sky130_fd_sc_hd__o2111ai_4 _39609_ (.A1(_16820_),
    .A2(_16823_),
    .B1(_16635_),
    .C1(_16631_),
    .D1(_16828_),
    .Y(_17030_));
 sky130_fd_sc_hd__nor2_1 _39610_ (.A(_17030_),
    .B(_16639_),
    .Y(_17031_));
 sky130_fd_sc_hd__and2_1 _39611_ (.A(_16242_),
    .B(_17031_),
    .X(_17032_));
 sky130_fd_sc_hd__or3_2 _39612_ (.A(_17023_),
    .B(_17029_),
    .C(_17032_),
    .X(_17033_));
 sky130_fd_sc_hd__o21ai_1 _39613_ (.A1(_17029_),
    .A2(_17032_),
    .B1(_17023_),
    .Y(_17034_));
 sky130_fd_sc_hd__and2_2 _39614_ (.A(_17033_),
    .B(_17034_),
    .X(_02671_));
 sky130_fd_sc_hd__nand2_2 _39615_ (.A(_17018_),
    .B(_17010_),
    .Y(_17035_));
 sky130_fd_sc_hd__a21oi_4 _39616_ (.A1(_16964_),
    .A2(_16969_),
    .B1(_16967_),
    .Y(_17036_));
 sky130_fd_sc_hd__a21oi_4 _39617_ (.A1(_16985_),
    .A2(_16970_),
    .B1(_17036_),
    .Y(_17037_));
 sky130_vsdinv _39618_ (.A(_16841_),
    .Y(_17038_));
 sky130_fd_sc_hd__o21a_2 _39619_ (.A1(_16509_),
    .A2(_16875_),
    .B1(_16873_),
    .X(_17039_));
 sky130_vsdinv _39620_ (.A(_17039_),
    .Y(_17040_));
 sky130_fd_sc_hd__a21o_1 _39621_ (.A1(_15813_),
    .A2(_16365_),
    .B1(_16839_),
    .X(_17041_));
 sky130_fd_sc_hd__nand2_1 _39622_ (.A(_17040_),
    .B(_17041_),
    .Y(_17042_));
 sky130_fd_sc_hd__nand2_1 _39623_ (.A(_17041_),
    .B(_16841_),
    .Y(_17043_));
 sky130_fd_sc_hd__nand2_1 _39624_ (.A(_17043_),
    .B(_17039_),
    .Y(_17044_));
 sky130_fd_sc_hd__o21ai_2 _39625_ (.A1(_17038_),
    .A2(_17042_),
    .B1(_17044_),
    .Y(_17045_));
 sky130_fd_sc_hd__nor2_2 _39626_ (.A(_15835_),
    .B(_17045_),
    .Y(_17046_));
 sky130_fd_sc_hd__and2_1 _39627_ (.A(_17045_),
    .B(_15834_),
    .X(_17047_));
 sky130_fd_sc_hd__or2_1 _39628_ (.A(_17046_),
    .B(_17047_),
    .X(_17048_));
 sky130_fd_sc_hd__a21oi_2 _39629_ (.A1(_16891_),
    .A2(_16894_),
    .B1(_17048_),
    .Y(_17049_));
 sky130_fd_sc_hd__nor2_4 _39630_ (.A(_17046_),
    .B(_17047_),
    .Y(_17050_));
 sky130_fd_sc_hd__nand2_2 _39631_ (.A(_16894_),
    .B(_16891_),
    .Y(_17051_));
 sky130_fd_sc_hd__nor2_4 _39632_ (.A(_17050_),
    .B(_17051_),
    .Y(_17052_));
 sky130_vsdinv _39633_ (.A(_16844_),
    .Y(_17053_));
 sky130_fd_sc_hd__and2_1 _39634_ (.A(_16846_),
    .B(_15835_),
    .X(_17054_));
 sky130_fd_sc_hd__nor2_4 _39635_ (.A(_17053_),
    .B(_17054_),
    .Y(_17055_));
 sky130_fd_sc_hd__o21a_1 _39636_ (.A1(_17049_),
    .A2(_17052_),
    .B1(_17055_),
    .X(_17056_));
 sky130_fd_sc_hd__nand2_4 _39637_ (.A(_17051_),
    .B(_17050_),
    .Y(_17057_));
 sky130_vsdinv _39638_ (.A(_17055_),
    .Y(_17058_));
 sky130_fd_sc_hd__nand2_1 _39639_ (.A(_17057_),
    .B(_17058_),
    .Y(_17059_));
 sky130_fd_sc_hd__nor2_4 _39640_ (.A(_17052_),
    .B(_17059_),
    .Y(_17060_));
 sky130_fd_sc_hd__nand2_2 _39641_ (.A(_11396_),
    .B(_11174_),
    .Y(_17061_));
 sky130_fd_sc_hd__nand2_2 _39642_ (.A(_12855_),
    .B(_10778_),
    .Y(_17062_));
 sky130_fd_sc_hd__or2_2 _39643_ (.A(_17061_),
    .B(_17062_),
    .X(_17063_));
 sky130_fd_sc_hd__nand2_2 _39644_ (.A(_17061_),
    .B(_17062_),
    .Y(_17064_));
 sky130_fd_sc_hd__nand2_2 _39645_ (.A(_11603_),
    .B(_19867_),
    .Y(_17065_));
 sky130_vsdinv _39646_ (.A(_17065_),
    .Y(_17066_));
 sky130_fd_sc_hd__a21o_1 _39647_ (.A1(_17063_),
    .A2(_17064_),
    .B1(_17066_),
    .X(_17067_));
 sky130_fd_sc_hd__nand3_4 _39648_ (.A(_17063_),
    .B(_17066_),
    .C(_17064_),
    .Y(_17068_));
 sky130_fd_sc_hd__o21bai_2 _39649_ (.A1(_16860_),
    .A2(_16864_),
    .B1_N(_16863_),
    .Y(_17069_));
 sky130_fd_sc_hd__a21o_1 _39650_ (.A1(_17067_),
    .A2(_17068_),
    .B1(_17069_),
    .X(_17070_));
 sky130_fd_sc_hd__nand3_4 _39651_ (.A(_17067_),
    .B(_17068_),
    .C(_17069_),
    .Y(_17071_));
 sky130_fd_sc_hd__a21oi_1 _39652_ (.A1(_17070_),
    .A2(_17071_),
    .B1(_16879_),
    .Y(_17072_));
 sky130_fd_sc_hd__and3_1 _39653_ (.A(_16879_),
    .B(_17070_),
    .C(_17071_),
    .X(_17073_));
 sky130_vsdinv _39654_ (.A(_16930_),
    .Y(_17074_));
 sky130_fd_sc_hd__a21oi_1 _39655_ (.A1(_16929_),
    .A2(_16931_),
    .B1(_17074_),
    .Y(_17075_));
 sky130_fd_sc_hd__o21ai_1 _39656_ (.A1(_17072_),
    .A2(_17073_),
    .B1(_17075_),
    .Y(_17076_));
 sky130_fd_sc_hd__a21o_1 _39657_ (.A1(_16929_),
    .A2(_16931_),
    .B1(_17074_),
    .X(_17077_));
 sky130_fd_sc_hd__a21o_1 _39658_ (.A1(_17070_),
    .A2(_17071_),
    .B1(_16879_),
    .X(_17078_));
 sky130_fd_sc_hd__nand3_4 _39659_ (.A(_16879_),
    .B(_17070_),
    .C(_17071_),
    .Y(_17079_));
 sky130_fd_sc_hd__nand3_4 _39660_ (.A(_17077_),
    .B(_17078_),
    .C(_17079_),
    .Y(_17080_));
 sky130_fd_sc_hd__nand2_1 _39661_ (.A(_17076_),
    .B(_17080_),
    .Y(_17081_));
 sky130_fd_sc_hd__a21oi_4 _39662_ (.A1(_16882_),
    .A2(_16879_),
    .B1(_16871_),
    .Y(_17082_));
 sky130_fd_sc_hd__and2_1 _39663_ (.A(_17081_),
    .B(_17082_),
    .X(_17083_));
 sky130_fd_sc_hd__a21oi_2 _39664_ (.A1(_17078_),
    .A2(_17079_),
    .B1(_17077_),
    .Y(_17084_));
 sky130_fd_sc_hd__nor2_1 _39665_ (.A(_17082_),
    .B(_17084_),
    .Y(_17085_));
 sky130_fd_sc_hd__nand2_2 _39666_ (.A(_17085_),
    .B(_17080_),
    .Y(_17086_));
 sky130_vsdinv _39667_ (.A(_17086_),
    .Y(_17087_));
 sky130_fd_sc_hd__nor2_2 _39668_ (.A(_10405_),
    .B(_12604_),
    .Y(_17088_));
 sky130_fd_sc_hd__and4_2 _39669_ (.A(_09733_),
    .B(_18695_),
    .C(_19830_),
    .D(_11085_),
    .X(_17089_));
 sky130_fd_sc_hd__o22a_2 _39670_ (.A1(_20109_),
    .A2(_15914_),
    .B1(_16103_),
    .B2(_12100_),
    .X(_17090_));
 sky130_fd_sc_hd__or3_4 _39671_ (.A(_17088_),
    .B(_17089_),
    .C(_17090_),
    .X(_17091_));
 sky130_fd_sc_hd__o21ai_4 _39672_ (.A1(_17089_),
    .A2(_17090_),
    .B1(_17088_),
    .Y(_17092_));
 sky130_fd_sc_hd__nor2_1 _39673_ (.A(_16896_),
    .B(_16897_),
    .Y(_17093_));
 sky130_fd_sc_hd__or2_4 _39674_ (.A(_16898_),
    .B(_17093_),
    .X(_17094_));
 sky130_fd_sc_hd__a21o_1 _39675_ (.A1(_17091_),
    .A2(_17092_),
    .B1(_17094_),
    .X(_17095_));
 sky130_fd_sc_hd__nand3_4 _39676_ (.A(_17094_),
    .B(_17092_),
    .C(_17091_),
    .Y(_17096_));
 sky130_fd_sc_hd__nor2_1 _39677_ (.A(_09321_),
    .B(_11941_),
    .Y(_17097_));
 sky130_fd_sc_hd__a22o_1 _39678_ (.A1(_19836_),
    .A2(_12304_),
    .B1(_15925_),
    .B2(_13451_),
    .X(_17098_));
 sky130_fd_sc_hd__o21a_1 _39679_ (.A1(_10988_),
    .A2(_12104_),
    .B1(_17098_),
    .X(_17099_));
 sky130_fd_sc_hd__or2_1 _39680_ (.A(_17097_),
    .B(_17099_),
    .X(_17100_));
 sky130_fd_sc_hd__nand2_1 _39681_ (.A(_17099_),
    .B(_17097_),
    .Y(_17101_));
 sky130_fd_sc_hd__and2_2 _39682_ (.A(_17100_),
    .B(_17101_),
    .X(_17102_));
 sky130_fd_sc_hd__a21bo_1 _39683_ (.A1(_17095_),
    .A2(_17096_),
    .B1_N(_17102_),
    .X(_17103_));
 sky130_fd_sc_hd__a21oi_4 _39684_ (.A1(_16904_),
    .A2(_16908_),
    .B1(_16914_),
    .Y(_17104_));
 sky130_fd_sc_hd__nand3b_2 _39685_ (.A_N(_17102_),
    .B(_17095_),
    .C(_17096_),
    .Y(_17105_));
 sky130_fd_sc_hd__nand3_4 _39686_ (.A(_17103_),
    .B(_17104_),
    .C(_17105_),
    .Y(_17106_));
 sky130_fd_sc_hd__a21o_1 _39687_ (.A1(_17095_),
    .A2(_17096_),
    .B1(_17102_),
    .X(_17107_));
 sky130_fd_sc_hd__nand3_2 _39688_ (.A(_17095_),
    .B(_17096_),
    .C(_17102_),
    .Y(_17108_));
 sky130_fd_sc_hd__nand3b_4 _39689_ (.A_N(_17104_),
    .B(_17107_),
    .C(_17108_),
    .Y(_17109_));
 sky130_fd_sc_hd__and4_4 _39690_ (.A(_19849_),
    .B(_19852_),
    .C(_20083_),
    .D(_20088_),
    .X(_17110_));
 sky130_fd_sc_hd__nand2_1 _39691_ (.A(_19855_),
    .B(_20080_),
    .Y(_17111_));
 sky130_fd_sc_hd__o22a_1 _39692_ (.A1(_16670_),
    .A2(_12297_),
    .B1(_15010_),
    .B2(_10763_),
    .X(_17112_));
 sky130_fd_sc_hd__or3_4 _39693_ (.A(_17110_),
    .B(_17111_),
    .C(_17112_),
    .X(_17113_));
 sky130_fd_sc_hd__o21ai_1 _39694_ (.A1(_17110_),
    .A2(_17112_),
    .B1(_17111_),
    .Y(_17114_));
 sky130_fd_sc_hd__nand2_1 _39695_ (.A(_17113_),
    .B(_17114_),
    .Y(_17115_));
 sky130_fd_sc_hd__o2bb2a_1 _39696_ (.A1_N(_16906_),
    .A2_N(_16905_),
    .B1(_16311_),
    .B2(_11737_),
    .X(_17116_));
 sky130_fd_sc_hd__nand2_2 _39697_ (.A(_17115_),
    .B(_17116_),
    .Y(_17117_));
 sky130_fd_sc_hd__nand3b_2 _39698_ (.A_N(_17116_),
    .B(_17113_),
    .C(_17114_),
    .Y(_17118_));
 sky130_fd_sc_hd__nand2_1 _39699_ (.A(_17117_),
    .B(_17118_),
    .Y(_17119_));
 sky130_vsdinv _39700_ (.A(_16927_),
    .Y(_17120_));
 sky130_fd_sc_hd__nor2_2 _39701_ (.A(_16923_),
    .B(_17120_),
    .Y(_17121_));
 sky130_fd_sc_hd__and2_1 _39702_ (.A(_17119_),
    .B(_17121_),
    .X(_17122_));
 sky130_fd_sc_hd__nor2_2 _39703_ (.A(_17121_),
    .B(_17119_),
    .Y(_17123_));
 sky130_fd_sc_hd__o2bb2ai_4 _39704_ (.A1_N(_17106_),
    .A2_N(_17109_),
    .B1(_17122_),
    .B2(_17123_),
    .Y(_17124_));
 sky130_fd_sc_hd__or2_2 _39705_ (.A(_16923_),
    .B(_17120_),
    .X(_17125_));
 sky130_fd_sc_hd__nand2_1 _39706_ (.A(_17119_),
    .B(_17125_),
    .Y(_17126_));
 sky130_fd_sc_hd__nand3_1 _39707_ (.A(_17117_),
    .B(_17121_),
    .C(_17118_),
    .Y(_17127_));
 sky130_fd_sc_hd__nand2_2 _39708_ (.A(_17126_),
    .B(_17127_),
    .Y(_17128_));
 sky130_fd_sc_hd__nand3_4 _39709_ (.A(_17109_),
    .B(_17106_),
    .C(_17128_),
    .Y(_17129_));
 sky130_fd_sc_hd__nand2_1 _39710_ (.A(_16919_),
    .B(_16935_),
    .Y(_17130_));
 sky130_fd_sc_hd__nand2_4 _39711_ (.A(_17130_),
    .B(_16913_),
    .Y(_17131_));
 sky130_fd_sc_hd__a21oi_4 _39712_ (.A1(_17124_),
    .A2(_17129_),
    .B1(_17131_),
    .Y(_17132_));
 sky130_fd_sc_hd__and3_1 _39713_ (.A(_17124_),
    .B(_17131_),
    .C(_17129_),
    .X(_17133_));
 sky130_fd_sc_hd__o22ai_4 _39714_ (.A1(_17083_),
    .A2(_17087_),
    .B1(_17132_),
    .B2(_17133_),
    .Y(_17134_));
 sky130_fd_sc_hd__nand2_1 _39715_ (.A(_17081_),
    .B(_17082_),
    .Y(_17135_));
 sky130_fd_sc_hd__nand2_2 _39716_ (.A(_17086_),
    .B(_17135_),
    .Y(_17136_));
 sky130_fd_sc_hd__a21o_1 _39717_ (.A1(_17124_),
    .A2(_17129_),
    .B1(_17131_),
    .X(_17137_));
 sky130_fd_sc_hd__nand3_4 _39718_ (.A(_17124_),
    .B(_17131_),
    .C(_17129_),
    .Y(_17138_));
 sky130_fd_sc_hd__nand3b_4 _39719_ (.A_N(_17136_),
    .B(_17137_),
    .C(_17138_),
    .Y(_17139_));
 sky130_fd_sc_hd__nand2_1 _39720_ (.A(_16887_),
    .B(_16891_),
    .Y(_17140_));
 sky130_fd_sc_hd__nand2_1 _39721_ (.A(_17140_),
    .B(_16948_),
    .Y(_17141_));
 sky130_fd_sc_hd__nand2_2 _39722_ (.A(_17141_),
    .B(_16894_),
    .Y(_17142_));
 sky130_fd_sc_hd__o21ai_4 _39723_ (.A1(_17142_),
    .A2(_16939_),
    .B1(_16947_),
    .Y(_17143_));
 sky130_fd_sc_hd__a21oi_4 _39724_ (.A1(_17134_),
    .A2(_17139_),
    .B1(_17143_),
    .Y(_17144_));
 sky130_fd_sc_hd__a21oi_1 _39725_ (.A1(_16944_),
    .A2(_16945_),
    .B1(_17142_),
    .Y(_17145_));
 sky130_fd_sc_hd__o211a_1 _39726_ (.A1(_16942_),
    .A2(_17145_),
    .B1(_17139_),
    .C1(_17134_),
    .X(_17146_));
 sky130_fd_sc_hd__o22ai_4 _39727_ (.A1(_17056_),
    .A2(_17060_),
    .B1(_17144_),
    .B2(_17146_),
    .Y(_17147_));
 sky130_fd_sc_hd__o21ai_2 _39728_ (.A1(_16968_),
    .A2(_16953_),
    .B1(_16961_),
    .Y(_17148_));
 sky130_fd_sc_hd__a21o_1 _39729_ (.A1(_17134_),
    .A2(_17139_),
    .B1(_17143_),
    .X(_17149_));
 sky130_fd_sc_hd__nor2_2 _39730_ (.A(_17060_),
    .B(_17056_),
    .Y(_17150_));
 sky130_fd_sc_hd__nand3_4 _39731_ (.A(_17134_),
    .B(_17143_),
    .C(_17139_),
    .Y(_17151_));
 sky130_fd_sc_hd__nand3_2 _39732_ (.A(_17149_),
    .B(_17150_),
    .C(_17151_),
    .Y(_17152_));
 sky130_fd_sc_hd__nand3_4 _39733_ (.A(_17147_),
    .B(_17148_),
    .C(_17152_),
    .Y(_17153_));
 sky130_fd_sc_hd__o21ai_2 _39734_ (.A1(_17144_),
    .A2(_17146_),
    .B1(_17150_),
    .Y(_17154_));
 sky130_fd_sc_hd__nand2_1 _39735_ (.A(_16961_),
    .B(_16968_),
    .Y(_17155_));
 sky130_fd_sc_hd__nand2_1 _39736_ (.A(_17155_),
    .B(_16957_),
    .Y(_17156_));
 sky130_fd_sc_hd__nand3b_4 _39737_ (.A_N(_17052_),
    .B(_17057_),
    .C(_17058_),
    .Y(_17157_));
 sky130_fd_sc_hd__o21ai_1 _39738_ (.A1(_17049_),
    .A2(_17052_),
    .B1(_17055_),
    .Y(_17158_));
 sky130_fd_sc_hd__nand2_2 _39739_ (.A(_17157_),
    .B(_17158_),
    .Y(_17159_));
 sky130_fd_sc_hd__nand3_2 _39740_ (.A(_17149_),
    .B(_17159_),
    .C(_17151_),
    .Y(_17160_));
 sky130_fd_sc_hd__nand3_4 _39741_ (.A(_17154_),
    .B(_17156_),
    .C(_17160_),
    .Y(_17161_));
 sky130_vsdinv _39742_ (.A(_16852_),
    .Y(_17162_));
 sky130_fd_sc_hd__o21ai_2 _39743_ (.A1(_17162_),
    .A2(_16859_),
    .B1(_16783_),
    .Y(_17163_));
 sky130_fd_sc_hd__a211o_1 _39744_ (.A1(_16855_),
    .A2(_16857_),
    .B1(_16256_),
    .C1(_17162_),
    .X(_17164_));
 sky130_fd_sc_hd__nand3_2 _39745_ (.A(_17163_),
    .B(_16982_),
    .C(_17164_),
    .Y(_17165_));
 sky130_vsdinv _39746_ (.A(_17165_),
    .Y(_17166_));
 sky130_fd_sc_hd__nand2_1 _39747_ (.A(_17163_),
    .B(_17164_),
    .Y(_17167_));
 sky130_fd_sc_hd__nand2_1 _39748_ (.A(_17167_),
    .B(_16787_),
    .Y(_17168_));
 sky130_vsdinv _39749_ (.A(_17168_),
    .Y(_17169_));
 sky130_fd_sc_hd__o2bb2ai_4 _39750_ (.A1_N(_17153_),
    .A2_N(_17161_),
    .B1(_17166_),
    .B2(_17169_),
    .Y(_17170_));
 sky130_fd_sc_hd__nand2_2 _39751_ (.A(_17168_),
    .B(_17165_),
    .Y(_17171_));
 sky130_fd_sc_hd__nand3b_4 _39752_ (.A_N(_17171_),
    .B(_17161_),
    .C(_17153_),
    .Y(_17172_));
 sky130_fd_sc_hd__nand3_4 _39753_ (.A(_17037_),
    .B(_17170_),
    .C(_17172_),
    .Y(_17173_));
 sky130_fd_sc_hd__a31oi_4 _39754_ (.A1(_16964_),
    .A2(_16967_),
    .A3(_16969_),
    .B1(_16984_),
    .Y(_17174_));
 sky130_fd_sc_hd__nand3_2 _39755_ (.A(_17161_),
    .B(_17153_),
    .C(_17171_),
    .Y(_17175_));
 sky130_fd_sc_hd__clkbuf_4 _39756_ (.A(_16982_),
    .X(_17176_));
 sky130_fd_sc_hd__nor2_1 _39757_ (.A(_17176_),
    .B(_17167_),
    .Y(_17177_));
 sky130_fd_sc_hd__and2_1 _39758_ (.A(_17167_),
    .B(_16992_),
    .X(_17178_));
 sky130_fd_sc_hd__o2bb2ai_2 _39759_ (.A1_N(_17153_),
    .A2_N(_17161_),
    .B1(_17177_),
    .B2(_17178_),
    .Y(_17179_));
 sky130_fd_sc_hd__o211ai_4 _39760_ (.A1(_17036_),
    .A2(_17174_),
    .B1(_17175_),
    .C1(_17179_),
    .Y(_17180_));
 sky130_fd_sc_hd__nand2_2 _39761_ (.A(_16978_),
    .B(_16972_),
    .Y(_17181_));
 sky130_fd_sc_hd__nor2_2 _39762_ (.A(net413),
    .B(_17181_),
    .Y(_17182_));
 sky130_vsdinv _39763_ (.A(_17181_),
    .Y(_17183_));
 sky130_fd_sc_hd__nor2_2 _39764_ (.A(_16426_),
    .B(_17183_),
    .Y(_17184_));
 sky130_fd_sc_hd__nor2_4 _39765_ (.A(_17182_),
    .B(_17184_),
    .Y(_17185_));
 sky130_fd_sc_hd__nand3_2 _39766_ (.A(_17173_),
    .B(_17180_),
    .C(_17185_),
    .Y(_17186_));
 sky130_fd_sc_hd__o2bb2ai_1 _39767_ (.A1_N(_17180_),
    .A2_N(_17173_),
    .B1(_17184_),
    .B2(_17182_),
    .Y(_17187_));
 sky130_fd_sc_hd__o2111ai_4 _39768_ (.A1(_16989_),
    .A2(_17000_),
    .B1(_16999_),
    .C1(_17186_),
    .D1(_17187_),
    .Y(_17188_));
 sky130_fd_sc_hd__o21ai_2 _39769_ (.A1(_17000_),
    .A2(_16989_),
    .B1(_16999_),
    .Y(_17189_));
 sky130_fd_sc_hd__nor2_2 _39770_ (.A(net413),
    .B(_17183_),
    .Y(_17190_));
 sky130_fd_sc_hd__clkbuf_2 _39771_ (.A(_17190_),
    .X(_17191_));
 sky130_fd_sc_hd__nor2_4 _39772_ (.A(_16426_),
    .B(_17181_),
    .Y(_17192_));
 sky130_fd_sc_hd__o2bb2ai_2 _39773_ (.A1_N(_17180_),
    .A2_N(_17173_),
    .B1(_17191_),
    .B2(_17192_),
    .Y(_17193_));
 sky130_fd_sc_hd__nor2_4 _39774_ (.A(_17192_),
    .B(_17190_),
    .Y(_17194_));
 sky130_fd_sc_hd__nand3_4 _39775_ (.A(_17173_),
    .B(_17180_),
    .C(_17194_),
    .Y(_17195_));
 sky130_fd_sc_hd__nand3_4 _39776_ (.A(_17189_),
    .B(_17193_),
    .C(_17195_),
    .Y(_17196_));
 sky130_fd_sc_hd__nand2_2 _39777_ (.A(_17188_),
    .B(_17196_),
    .Y(_17197_));
 sky130_vsdinv _39778_ (.A(_17003_),
    .Y(_17198_));
 sky130_fd_sc_hd__nand2_2 _39779_ (.A(_17197_),
    .B(_17198_),
    .Y(_17199_));
 sky130_fd_sc_hd__nand3_4 _39780_ (.A(_17188_),
    .B(_17196_),
    .C(_17003_),
    .Y(_17200_));
 sky130_fd_sc_hd__nand3_4 _39781_ (.A(_17035_),
    .B(_17199_),
    .C(_17200_),
    .Y(_17201_));
 sky130_fd_sc_hd__nand2_1 _39782_ (.A(_17197_),
    .B(_17003_),
    .Y(_17202_));
 sky130_fd_sc_hd__a21boi_2 _39783_ (.A1(_17002_),
    .A2(_17011_),
    .B1_N(_17010_),
    .Y(_17203_));
 sky130_fd_sc_hd__nand3_2 _39784_ (.A(_17188_),
    .B(_17196_),
    .C(_17198_),
    .Y(_17204_));
 sky130_fd_sc_hd__nand3_4 _39785_ (.A(_17202_),
    .B(_17203_),
    .C(_17204_),
    .Y(_17205_));
 sky130_fd_sc_hd__nand2_2 _39786_ (.A(_17201_),
    .B(_17205_),
    .Y(_17206_));
 sky130_fd_sc_hd__nand2_2 _39787_ (.A(_17034_),
    .B(_17022_),
    .Y(_17207_));
 sky130_fd_sc_hd__xnor2_4 _39788_ (.A(_17206_),
    .B(_17207_),
    .Y(_02672_));
 sky130_vsdinv _39789_ (.A(_17200_),
    .Y(_17208_));
 sky130_fd_sc_hd__a31oi_2 _39790_ (.A1(_16832_),
    .A2(_16997_),
    .A3(_17001_),
    .B1(_17020_),
    .Y(_17209_));
 sky130_fd_sc_hd__o2bb2ai_2 _39791_ (.A1_N(_17198_),
    .A2_N(_17197_),
    .B1(_17017_),
    .B2(_17209_),
    .Y(_17210_));
 sky130_fd_sc_hd__o2111a_1 _39792_ (.A1(_17208_),
    .A2(_17210_),
    .B1(_17022_),
    .C1(_17205_),
    .D1(_17016_),
    .X(_17211_));
 sky130_fd_sc_hd__o21ai_2 _39793_ (.A1(_17029_),
    .A2(_17032_),
    .B1(_17211_),
    .Y(_17212_));
 sky130_fd_sc_hd__a21oi_2 _39794_ (.A1(_17199_),
    .A2(_17200_),
    .B1(_17035_),
    .Y(_17213_));
 sky130_fd_sc_hd__a21oi_4 _39795_ (.A1(_17022_),
    .A2(_17201_),
    .B1(_17213_),
    .Y(_17214_));
 sky130_vsdinv _39796_ (.A(_17214_),
    .Y(_17215_));
 sky130_fd_sc_hd__a21oi_4 _39797_ (.A1(_17170_),
    .A2(_17172_),
    .B1(_17037_),
    .Y(_17216_));
 sky130_fd_sc_hd__a31oi_4 _39798_ (.A1(_17037_),
    .A2(_17170_),
    .A3(_17172_),
    .B1(_17185_),
    .Y(_17217_));
 sky130_vsdinv _39799_ (.A(_17118_),
    .Y(_17218_));
 sky130_fd_sc_hd__a21o_1 _39800_ (.A1(_17125_),
    .A2(_17117_),
    .B1(_17218_),
    .X(_17219_));
 sky130_fd_sc_hd__nand2_2 _39801_ (.A(_19860_),
    .B(_20070_),
    .Y(_17220_));
 sky130_fd_sc_hd__nand2_2 _39802_ (.A(_11603_),
    .B(_19864_),
    .Y(_17221_));
 sky130_fd_sc_hd__xor2_1 _39803_ (.A(_17220_),
    .B(_17221_),
    .X(_17222_));
 sky130_fd_sc_hd__or2_1 _39804_ (.A(_17066_),
    .B(_17222_),
    .X(_17223_));
 sky130_fd_sc_hd__nand2_1 _39805_ (.A(_17222_),
    .B(_17066_),
    .Y(_17224_));
 sky130_fd_sc_hd__nand2_1 _39806_ (.A(_17068_),
    .B(_17063_),
    .Y(_17225_));
 sky130_vsdinv _39807_ (.A(_17225_),
    .Y(_17226_));
 sky130_fd_sc_hd__a21o_1 _39808_ (.A1(_17223_),
    .A2(_17224_),
    .B1(_17226_),
    .X(_17227_));
 sky130_fd_sc_hd__xor2_1 _39809_ (.A(_17065_),
    .B(_17221_),
    .X(_17228_));
 sky130_fd_sc_hd__or2_2 _39810_ (.A(_17220_),
    .B(_17228_),
    .X(_17229_));
 sky130_fd_sc_hd__nand2_1 _39811_ (.A(_17228_),
    .B(_17220_),
    .Y(_17230_));
 sky130_fd_sc_hd__a21o_1 _39812_ (.A1(_17229_),
    .A2(_17230_),
    .B1(_17225_),
    .X(_17231_));
 sky130_fd_sc_hd__nand3_4 _39813_ (.A(_17227_),
    .B(_17231_),
    .C(_16885_),
    .Y(_17232_));
 sky130_fd_sc_hd__a21o_1 _39814_ (.A1(_17229_),
    .A2(_17230_),
    .B1(_17226_),
    .X(_17233_));
 sky130_fd_sc_hd__nand3_2 _39815_ (.A(_17229_),
    .B(_17226_),
    .C(_17230_),
    .Y(_17234_));
 sky130_fd_sc_hd__nand3_4 _39816_ (.A(_17233_),
    .B(_16878_),
    .C(_17234_),
    .Y(_17235_));
 sky130_fd_sc_hd__nand3_4 _39817_ (.A(_17219_),
    .B(_17232_),
    .C(_17235_),
    .Y(_17236_));
 sky130_fd_sc_hd__nand2_1 _39818_ (.A(_17232_),
    .B(_17235_),
    .Y(_17237_));
 sky130_fd_sc_hd__a21oi_2 _39819_ (.A1(_17125_),
    .A2(_17117_),
    .B1(_17218_),
    .Y(_17238_));
 sky130_fd_sc_hd__nand2_4 _39820_ (.A(_17237_),
    .B(_17238_),
    .Y(_17239_));
 sky130_fd_sc_hd__nand2_2 _39821_ (.A(_17079_),
    .B(_17071_),
    .Y(_17240_));
 sky130_fd_sc_hd__a21oi_4 _39822_ (.A1(_17236_),
    .A2(_17239_),
    .B1(_17240_),
    .Y(_17241_));
 sky130_fd_sc_hd__nand2_4 _39823_ (.A(_17239_),
    .B(_17240_),
    .Y(_17242_));
 sky130_vsdinv _39824_ (.A(_17236_),
    .Y(_17243_));
 sky130_fd_sc_hd__nor2_4 _39825_ (.A(_17242_),
    .B(_17243_),
    .Y(_17244_));
 sky130_fd_sc_hd__nand2_2 _39826_ (.A(_16107_),
    .B(_20099_),
    .Y(_17245_));
 sky130_fd_sc_hd__and4_2 _39827_ (.A(_08038_),
    .B(_13837_),
    .C(_19830_),
    .D(_12303_),
    .X(_17246_));
 sky130_fd_sc_hd__o22a_2 _39828_ (.A1(_11085_),
    .A2(_11275_),
    .B1(_16102_),
    .B2(_12604_),
    .X(_17247_));
 sky130_fd_sc_hd__nor2_4 _39829_ (.A(_17246_),
    .B(_17247_),
    .Y(_17248_));
 sky130_fd_sc_hd__or2_4 _39830_ (.A(_17245_),
    .B(_17248_),
    .X(_17249_));
 sky130_fd_sc_hd__nand2_4 _39831_ (.A(_17248_),
    .B(_17245_),
    .Y(_17250_));
 sky130_vsdinv _39832_ (.A(_17089_),
    .Y(_17251_));
 sky130_fd_sc_hd__o31a_2 _39833_ (.A1(_10405_),
    .A2(_12604_),
    .A3(_17090_),
    .B1(_17251_),
    .X(_17252_));
 sky130_fd_sc_hd__a21oi_4 _39834_ (.A1(_17249_),
    .A2(_17250_),
    .B1(_17252_),
    .Y(_17253_));
 sky130_fd_sc_hd__nand3_4 _39835_ (.A(_17249_),
    .B(_17250_),
    .C(_17252_),
    .Y(_17254_));
 sky130_vsdinv _39836_ (.A(_17254_),
    .Y(_17255_));
 sky130_fd_sc_hd__nand2_4 _39837_ (.A(_15897_),
    .B(_20088_),
    .Y(_17256_));
 sky130_fd_sc_hd__o22a_1 _39838_ (.A1(_16094_),
    .A2(_11557_),
    .B1(_16095_),
    .B2(_10781_),
    .X(_17257_));
 sky130_fd_sc_hd__a31o_1 _39839_ (.A1(_20092_),
    .A2(_20095_),
    .A3(_16092_),
    .B1(_17257_),
    .X(_17258_));
 sky130_fd_sc_hd__nor2_2 _39840_ (.A(_17256_),
    .B(_17258_),
    .Y(_17259_));
 sky130_fd_sc_hd__nand2_1 _39841_ (.A(_17258_),
    .B(_17256_),
    .Y(_17260_));
 sky130_fd_sc_hd__or2b_2 _39842_ (.A(_17259_),
    .B_N(_17260_),
    .X(_17261_));
 sky130_fd_sc_hd__o21ai_2 _39843_ (.A1(_17253_),
    .A2(_17255_),
    .B1(_17261_),
    .Y(_17262_));
 sky130_fd_sc_hd__a21oi_4 _39844_ (.A1(_17091_),
    .A2(_17092_),
    .B1(_17094_),
    .Y(_17263_));
 sky130_fd_sc_hd__a21o_1 _39845_ (.A1(_17102_),
    .A2(_17096_),
    .B1(_17263_),
    .X(_17264_));
 sky130_fd_sc_hd__nand2_1 _39846_ (.A(_17249_),
    .B(_17250_),
    .Y(_17265_));
 sky130_vsdinv _39847_ (.A(_17252_),
    .Y(_17266_));
 sky130_fd_sc_hd__nand2_2 _39848_ (.A(_17265_),
    .B(_17266_),
    .Y(_17267_));
 sky130_fd_sc_hd__and2_1 _39849_ (.A(_17258_),
    .B(_17256_),
    .X(_17268_));
 sky130_fd_sc_hd__nor2_4 _39850_ (.A(_17259_),
    .B(_17268_),
    .Y(_17269_));
 sky130_fd_sc_hd__nand3_4 _39851_ (.A(_17267_),
    .B(_17254_),
    .C(_17269_),
    .Y(_17270_));
 sky130_fd_sc_hd__nand3_4 _39852_ (.A(_17262_),
    .B(_17264_),
    .C(_17270_),
    .Y(_17271_));
 sky130_fd_sc_hd__o21ai_2 _39853_ (.A1(_17253_),
    .A2(_17255_),
    .B1(_17269_),
    .Y(_17272_));
 sky130_fd_sc_hd__a21oi_4 _39854_ (.A1(_17102_),
    .A2(_17096_),
    .B1(_17263_),
    .Y(_17273_));
 sky130_fd_sc_hd__nand3_4 _39855_ (.A(_17267_),
    .B(_17261_),
    .C(_17254_),
    .Y(_17274_));
 sky130_fd_sc_hd__nand3_4 _39856_ (.A(_17272_),
    .B(_17273_),
    .C(_17274_),
    .Y(_17275_));
 sky130_fd_sc_hd__nor2_4 _39857_ (.A(_08615_),
    .B(_16059_),
    .Y(_17276_));
 sky130_fd_sc_hd__nand2_4 _39858_ (.A(_19849_),
    .B(_11165_),
    .Y(_17277_));
 sky130_fd_sc_hd__nand2_4 _39859_ (.A(_19852_),
    .B(_13647_),
    .Y(_17278_));
 sky130_fd_sc_hd__xor2_4 _39860_ (.A(_17277_),
    .B(_17278_),
    .X(_17279_));
 sky130_fd_sc_hd__or2_4 _39861_ (.A(_17276_),
    .B(_17279_),
    .X(_17280_));
 sky130_fd_sc_hd__nand2_4 _39862_ (.A(_17279_),
    .B(_17276_),
    .Y(_17281_));
 sky130_fd_sc_hd__o21ai_4 _39863_ (.A1(_16327_),
    .A2(_12104_),
    .B1(_17101_),
    .Y(_17282_));
 sky130_fd_sc_hd__a21o_1 _39864_ (.A1(_17280_),
    .A2(_17281_),
    .B1(_17282_),
    .X(_17283_));
 sky130_fd_sc_hd__nand3_4 _39865_ (.A(_17280_),
    .B(_17282_),
    .C(_17281_),
    .Y(_17284_));
 sky130_fd_sc_hd__nand2_1 _39866_ (.A(_17283_),
    .B(_17284_),
    .Y(_17285_));
 sky130_vsdinv _39867_ (.A(_17113_),
    .Y(_17286_));
 sky130_fd_sc_hd__nor2_8 _39868_ (.A(_17110_),
    .B(_17286_),
    .Y(_17287_));
 sky130_fd_sc_hd__and2_1 _39869_ (.A(_17285_),
    .B(_17287_),
    .X(_17288_));
 sky130_fd_sc_hd__nor2_2 _39870_ (.A(_17287_),
    .B(_17285_),
    .Y(_17289_));
 sky130_fd_sc_hd__o2bb2ai_4 _39871_ (.A1_N(_17271_),
    .A2_N(_17275_),
    .B1(_17288_),
    .B2(_17289_),
    .Y(_17290_));
 sky130_fd_sc_hd__o21ai_1 _39872_ (.A1(_17110_),
    .A2(_17286_),
    .B1(_17285_),
    .Y(_17291_));
 sky130_fd_sc_hd__nand3_2 _39873_ (.A(_17287_),
    .B(_17283_),
    .C(_17284_),
    .Y(_17292_));
 sky130_fd_sc_hd__nand2_2 _39874_ (.A(_17291_),
    .B(_17292_),
    .Y(_17293_));
 sky130_fd_sc_hd__nand3_4 _39875_ (.A(_17271_),
    .B(_17275_),
    .C(_17293_),
    .Y(_17294_));
 sky130_fd_sc_hd__nand2_1 _39876_ (.A(_17106_),
    .B(_17128_),
    .Y(_17295_));
 sky130_fd_sc_hd__nand2_4 _39877_ (.A(_17295_),
    .B(_17109_),
    .Y(_17296_));
 sky130_fd_sc_hd__a21oi_4 _39878_ (.A1(_17290_),
    .A2(_17294_),
    .B1(_17296_),
    .Y(_17297_));
 sky130_fd_sc_hd__and3_2 _39879_ (.A(_17290_),
    .B(_17296_),
    .C(_17294_),
    .X(_17298_));
 sky130_fd_sc_hd__o22ai_4 _39880_ (.A1(_17241_),
    .A2(_17244_),
    .B1(_17297_),
    .B2(_17298_),
    .Y(_17299_));
 sky130_fd_sc_hd__nand2_1 _39881_ (.A(_17290_),
    .B(_17294_),
    .Y(_17300_));
 sky130_vsdinv _39882_ (.A(_17296_),
    .Y(_17301_));
 sky130_fd_sc_hd__nand2_2 _39883_ (.A(_17300_),
    .B(_17301_),
    .Y(_17302_));
 sky130_fd_sc_hd__nor2_4 _39884_ (.A(_17241_),
    .B(_17244_),
    .Y(_17303_));
 sky130_fd_sc_hd__nand3_4 _39885_ (.A(_17290_),
    .B(_17296_),
    .C(_17294_),
    .Y(_17304_));
 sky130_fd_sc_hd__nand3_4 _39886_ (.A(_17302_),
    .B(_17303_),
    .C(_17304_),
    .Y(_17305_));
 sky130_fd_sc_hd__o21ai_2 _39887_ (.A1(_17136_),
    .A2(_17132_),
    .B1(_17138_),
    .Y(_17306_));
 sky130_fd_sc_hd__nand3_4 _39888_ (.A(_17299_),
    .B(_17305_),
    .C(_17306_),
    .Y(_17307_));
 sky130_fd_sc_hd__o21ai_2 _39889_ (.A1(_17297_),
    .A2(_17298_),
    .B1(_17303_),
    .Y(_17308_));
 sky130_fd_sc_hd__o21a_1 _39890_ (.A1(_17136_),
    .A2(_17132_),
    .B1(_17138_),
    .X(_17309_));
 sky130_fd_sc_hd__a21o_1 _39891_ (.A1(_17236_),
    .A2(_17239_),
    .B1(_17240_),
    .X(_17310_));
 sky130_fd_sc_hd__o21ai_4 _39892_ (.A1(_17243_),
    .A2(_17242_),
    .B1(_17310_),
    .Y(_17311_));
 sky130_fd_sc_hd__nand3_2 _39893_ (.A(_17302_),
    .B(_17311_),
    .C(_17304_),
    .Y(_17312_));
 sky130_fd_sc_hd__nand3_4 _39894_ (.A(_17308_),
    .B(_17309_),
    .C(_17312_),
    .Y(_17313_));
 sky130_fd_sc_hd__or2_4 _39895_ (.A(_16840_),
    .B(_17040_),
    .X(_17314_));
 sky130_fd_sc_hd__nor2_8 _39896_ (.A(_16841_),
    .B(_17039_),
    .Y(_17315_));
 sky130_vsdinv _39897_ (.A(_17315_),
    .Y(_17316_));
 sky130_fd_sc_hd__a21oi_4 _39898_ (.A1(_17314_),
    .A2(_17316_),
    .B1(_15834_),
    .Y(_17317_));
 sky130_fd_sc_hd__and3_2 _39899_ (.A(_17314_),
    .B(_15834_),
    .C(_17316_),
    .X(_17318_));
 sky130_fd_sc_hd__nor2_4 _39900_ (.A(_17317_),
    .B(_17318_),
    .Y(_17319_));
 sky130_fd_sc_hd__inv_4 _39901_ (.A(_17319_),
    .Y(_17320_));
 sky130_fd_sc_hd__nand3_4 _39902_ (.A(_17320_),
    .B(_17086_),
    .C(_17080_),
    .Y(_17321_));
 sky130_fd_sc_hd__o21ai_2 _39903_ (.A1(_17082_),
    .A2(_17084_),
    .B1(_17080_),
    .Y(_17322_));
 sky130_fd_sc_hd__buf_2 _39904_ (.A(_17319_),
    .X(_17323_));
 sky130_fd_sc_hd__nand2_2 _39905_ (.A(_17322_),
    .B(_17323_),
    .Y(_17324_));
 sky130_fd_sc_hd__nor2_2 _39906_ (.A(_17315_),
    .B(_17047_),
    .Y(_17325_));
 sky130_vsdinv _39907_ (.A(_17325_),
    .Y(_17326_));
 sky130_fd_sc_hd__a21oi_4 _39908_ (.A1(_17321_),
    .A2(_17324_),
    .B1(_17326_),
    .Y(_17327_));
 sky130_fd_sc_hd__and3_1 _39909_ (.A(_17321_),
    .B(_17326_),
    .C(_17324_),
    .X(_17328_));
 sky130_fd_sc_hd__o2bb2ai_4 _39910_ (.A1_N(_17307_),
    .A2_N(_17313_),
    .B1(_17327_),
    .B2(_17328_),
    .Y(_17329_));
 sky130_fd_sc_hd__and2_1 _39911_ (.A(_17324_),
    .B(_17326_),
    .X(_17330_));
 sky130_fd_sc_hd__a21oi_4 _39912_ (.A1(_17330_),
    .A2(_17321_),
    .B1(_17327_),
    .Y(_17331_));
 sky130_fd_sc_hd__nand3_4 _39913_ (.A(_17313_),
    .B(_17307_),
    .C(_17331_),
    .Y(_17332_));
 sky130_fd_sc_hd__o21ai_4 _39914_ (.A1(_17159_),
    .A2(_17144_),
    .B1(_17151_),
    .Y(_17333_));
 sky130_fd_sc_hd__a21oi_4 _39915_ (.A1(_17329_),
    .A2(_17332_),
    .B1(_17333_),
    .Y(_17334_));
 sky130_fd_sc_hd__and2_1 _39916_ (.A(_17134_),
    .B(_17139_),
    .X(_17335_));
 sky130_fd_sc_hd__nand2_1 _39917_ (.A(_17159_),
    .B(_17151_),
    .Y(_17336_));
 sky130_fd_sc_hd__o2111a_2 _39918_ (.A1(_17143_),
    .A2(_17335_),
    .B1(_17336_),
    .C1(_17332_),
    .D1(_17329_),
    .X(_17337_));
 sky130_fd_sc_hd__nand3_4 _39919_ (.A(_17157_),
    .B(_16258_),
    .C(_17057_),
    .Y(_17338_));
 sky130_fd_sc_hd__o21ai_1 _39920_ (.A1(_17055_),
    .A2(_17052_),
    .B1(_17057_),
    .Y(_17339_));
 sky130_fd_sc_hd__nand2_2 _39921_ (.A(_17339_),
    .B(_16783_),
    .Y(_17340_));
 sky130_fd_sc_hd__nand2_1 _39922_ (.A(_17338_),
    .B(_17340_),
    .Y(_17341_));
 sky130_fd_sc_hd__nand2_1 _39923_ (.A(_17341_),
    .B(_16982_),
    .Y(_17342_));
 sky130_fd_sc_hd__nand3_2 _39924_ (.A(_17338_),
    .B(_17340_),
    .C(_16787_),
    .Y(_17343_));
 sky130_fd_sc_hd__nand2_4 _39925_ (.A(_17342_),
    .B(_17343_),
    .Y(_17344_));
 sky130_fd_sc_hd__o21ai_2 _39926_ (.A1(_17334_),
    .A2(_17337_),
    .B1(_17344_),
    .Y(_17345_));
 sky130_fd_sc_hd__nand2_1 _39927_ (.A(_17161_),
    .B(_17171_),
    .Y(_17346_));
 sky130_fd_sc_hd__nand2_1 _39928_ (.A(_17346_),
    .B(_17153_),
    .Y(_17347_));
 sky130_fd_sc_hd__nand2_1 _39929_ (.A(_17329_),
    .B(_17332_),
    .Y(_17348_));
 sky130_fd_sc_hd__nand2_1 _39930_ (.A(_17336_),
    .B(_17149_),
    .Y(_17349_));
 sky130_fd_sc_hd__nand2_1 _39931_ (.A(_17348_),
    .B(_17349_),
    .Y(_17350_));
 sky130_fd_sc_hd__nand3_4 _39932_ (.A(_17333_),
    .B(_17329_),
    .C(_17332_),
    .Y(_17351_));
 sky130_fd_sc_hd__nand3b_2 _39933_ (.A_N(_17344_),
    .B(_17350_),
    .C(_17351_),
    .Y(_17352_));
 sky130_fd_sc_hd__nand3_4 _39934_ (.A(_17345_),
    .B(_17347_),
    .C(_17352_),
    .Y(_17353_));
 sky130_fd_sc_hd__nand2_1 _39935_ (.A(_17341_),
    .B(_16975_),
    .Y(_17354_));
 sky130_vsdinv _39936_ (.A(_17354_),
    .Y(_17355_));
 sky130_fd_sc_hd__nand3_1 _39937_ (.A(_17338_),
    .B(_17340_),
    .C(_16992_),
    .Y(_17356_));
 sky130_vsdinv _39938_ (.A(_17356_),
    .Y(_17357_));
 sky130_fd_sc_hd__o22ai_4 _39939_ (.A1(_17355_),
    .A2(_17357_),
    .B1(_17334_),
    .B2(_17337_),
    .Y(_17358_));
 sky130_fd_sc_hd__a21boi_2 _39940_ (.A1(_17161_),
    .A2(_17171_),
    .B1_N(_17153_),
    .Y(_17359_));
 sky130_fd_sc_hd__nand3_2 _39941_ (.A(_17350_),
    .B(_17351_),
    .C(_17344_),
    .Y(_17360_));
 sky130_fd_sc_hd__nand3_4 _39942_ (.A(_17358_),
    .B(_17359_),
    .C(_17360_),
    .Y(_17361_));
 sky130_fd_sc_hd__nand2_1 _39943_ (.A(_17164_),
    .B(_16592_),
    .Y(_17362_));
 sky130_fd_sc_hd__nand2_2 _39944_ (.A(_17362_),
    .B(_17163_),
    .Y(_17363_));
 sky130_fd_sc_hd__nor2_4 _39945_ (.A(_16423_),
    .B(_17363_),
    .Y(_17364_));
 sky130_vsdinv _39946_ (.A(_17363_),
    .Y(_17365_));
 sky130_fd_sc_hd__nor2_8 _39947_ (.A(_15754_),
    .B(_17365_),
    .Y(_17366_));
 sky130_fd_sc_hd__nor2_4 _39948_ (.A(_17364_),
    .B(_17366_),
    .Y(_17367_));
 sky130_fd_sc_hd__nand3_2 _39949_ (.A(_17353_),
    .B(_17361_),
    .C(_17367_),
    .Y(_17368_));
 sky130_fd_sc_hd__o2bb2ai_2 _39950_ (.A1_N(_17361_),
    .A2_N(_17353_),
    .B1(_17366_),
    .B2(_17364_),
    .Y(_17369_));
 sky130_fd_sc_hd__o211ai_4 _39951_ (.A1(_17216_),
    .A2(_17217_),
    .B1(_17368_),
    .C1(_17369_),
    .Y(_17370_));
 sky130_fd_sc_hd__nor2_1 _39952_ (.A(net412),
    .B(_17363_),
    .Y(_17371_));
 sky130_fd_sc_hd__nor2_1 _39953_ (.A(_17004_),
    .B(_17365_),
    .Y(_17372_));
 sky130_fd_sc_hd__o2bb2ai_2 _39954_ (.A1_N(_17361_),
    .A2_N(_17353_),
    .B1(_17371_),
    .B2(_17372_),
    .Y(_17373_));
 sky130_fd_sc_hd__a21oi_2 _39955_ (.A1(_17173_),
    .A2(_17194_),
    .B1(_17216_),
    .Y(_17374_));
 sky130_fd_sc_hd__nand3b_2 _39956_ (.A_N(_17367_),
    .B(_17353_),
    .C(_17361_),
    .Y(_17375_));
 sky130_fd_sc_hd__nand3_4 _39957_ (.A(_17373_),
    .B(_17374_),
    .C(_17375_),
    .Y(_17376_));
 sky130_fd_sc_hd__a21oi_1 _39958_ (.A1(_17370_),
    .A2(_17376_),
    .B1(_17191_),
    .Y(_17377_));
 sky130_fd_sc_hd__and3_1 _39959_ (.A(_17370_),
    .B(_17376_),
    .C(_17191_),
    .X(_17378_));
 sky130_fd_sc_hd__a21oi_1 _39960_ (.A1(_17193_),
    .A2(_17195_),
    .B1(_17189_),
    .Y(_17379_));
 sky130_fd_sc_hd__o21ai_2 _39961_ (.A1(_17198_),
    .A2(_17379_),
    .B1(_17196_),
    .Y(_17380_));
 sky130_fd_sc_hd__o21bai_2 _39962_ (.A1(_17377_),
    .A2(_17378_),
    .B1_N(_17380_),
    .Y(_17381_));
 sky130_fd_sc_hd__a21o_1 _39963_ (.A1(_17370_),
    .A2(_17376_),
    .B1(_17191_),
    .X(_17382_));
 sky130_fd_sc_hd__nand3_2 _39964_ (.A(_17370_),
    .B(_17376_),
    .C(_17191_),
    .Y(_17383_));
 sky130_fd_sc_hd__nand3_4 _39965_ (.A(_17382_),
    .B(_17380_),
    .C(_17383_),
    .Y(_17384_));
 sky130_fd_sc_hd__and2_2 _39966_ (.A(_17381_),
    .B(_17384_),
    .X(_17385_));
 sky130_fd_sc_hd__a21boi_4 _39967_ (.A1(_17212_),
    .A2(_17215_),
    .B1_N(_17385_),
    .Y(_17386_));
 sky130_fd_sc_hd__and3b_1 _39968_ (.A_N(_17385_),
    .B(_17212_),
    .C(_17215_),
    .X(_17387_));
 sky130_fd_sc_hd__nor2_4 _39969_ (.A(_17386_),
    .B(_17387_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand3_4 _39970_ (.A(_17320_),
    .B(_17236_),
    .C(_17242_),
    .Y(_17388_));
 sky130_fd_sc_hd__nand2_1 _39971_ (.A(_17242_),
    .B(_17236_),
    .Y(_17389_));
 sky130_fd_sc_hd__nand2_2 _39972_ (.A(_17389_),
    .B(_17323_),
    .Y(_17390_));
 sky130_fd_sc_hd__nor2_4 _39973_ (.A(_17315_),
    .B(_17318_),
    .Y(_17391_));
 sky130_vsdinv _39974_ (.A(_17391_),
    .Y(_17392_));
 sky130_fd_sc_hd__clkbuf_4 _39975_ (.A(_17392_),
    .X(_17393_));
 sky130_fd_sc_hd__a21oi_4 _39976_ (.A1(_17388_),
    .A2(_17390_),
    .B1(_17393_),
    .Y(_17394_));
 sky130_fd_sc_hd__and3_2 _39977_ (.A(_17388_),
    .B(_17390_),
    .C(_17392_),
    .X(_17395_));
 sky130_fd_sc_hd__a21oi_4 _39978_ (.A1(_17280_),
    .A2(_17281_),
    .B1(_17282_),
    .Y(_17396_));
 sky130_fd_sc_hd__o21ai_1 _39979_ (.A1(_19864_),
    .A2(_19868_),
    .B1(_19860_),
    .Y(_17397_));
 sky130_fd_sc_hd__a21oi_1 _39980_ (.A1(_19864_),
    .A2(_19868_),
    .B1(_16147_),
    .Y(_17398_));
 sky130_fd_sc_hd__o31a_2 _39981_ (.A1(_19860_),
    .A2(_19864_),
    .A3(_19868_),
    .B1(_18688_),
    .X(_17399_));
 sky130_fd_sc_hd__o21ai_2 _39982_ (.A1(_17397_),
    .A2(_17398_),
    .B1(_17399_),
    .Y(_17400_));
 sky130_fd_sc_hd__nor2_1 _39983_ (.A(_17400_),
    .B(_16885_),
    .Y(_17401_));
 sky130_fd_sc_hd__nand2_1 _39984_ (.A(_16885_),
    .B(_17400_),
    .Y(_17402_));
 sky130_fd_sc_hd__and2b_1 _39985_ (.A_N(_17401_),
    .B(_17402_),
    .X(_17403_));
 sky130_fd_sc_hd__o211ai_4 _39986_ (.A1(_17287_),
    .A2(_17396_),
    .B1(_17284_),
    .C1(_17403_),
    .Y(_17404_));
 sky130_fd_sc_hd__or2b_1 _39987_ (.A(_17401_),
    .B_N(_17402_),
    .X(_17405_));
 sky130_fd_sc_hd__o21ai_2 _39988_ (.A1(_17396_),
    .A2(_17287_),
    .B1(_17284_),
    .Y(_17406_));
 sky130_fd_sc_hd__nand2_2 _39989_ (.A(_17405_),
    .B(_17406_),
    .Y(_17407_));
 sky130_fd_sc_hd__and2_2 _39990_ (.A(_17235_),
    .B(_17233_),
    .X(_17408_));
 sky130_fd_sc_hd__and3_1 _39991_ (.A(_17404_),
    .B(_17407_),
    .C(_17408_),
    .X(_17409_));
 sky130_fd_sc_hd__a21oi_4 _39992_ (.A1(_17404_),
    .A2(_17407_),
    .B1(_17408_),
    .Y(_17410_));
 sky130_fd_sc_hd__nand2_1 _39993_ (.A(_19849_),
    .B(_13647_),
    .Y(_17411_));
 sky130_fd_sc_hd__nor2_2 _39994_ (.A(_15009_),
    .B(_10772_),
    .Y(_17412_));
 sky130_fd_sc_hd__or2_2 _39995_ (.A(_17411_),
    .B(_17412_),
    .X(_17413_));
 sky130_fd_sc_hd__nand2_2 _39996_ (.A(_17412_),
    .B(_17411_),
    .Y(_17414_));
 sky130_fd_sc_hd__nand2_2 _39997_ (.A(_19856_),
    .B(_20071_),
    .Y(_17415_));
 sky130_fd_sc_hd__a21o_2 _39998_ (.A1(_17413_),
    .A2(_17414_),
    .B1(_17415_),
    .X(_17416_));
 sky130_fd_sc_hd__nand3_4 _39999_ (.A(_17413_),
    .B(_17415_),
    .C(_17414_),
    .Y(_17417_));
 sky130_fd_sc_hd__o32ai_4 _40000_ (.A1(_11941_),
    .A2(_11563_),
    .A3(_16327_),
    .B1(_17256_),
    .B2(_17257_),
    .Y(_17418_));
 sky130_fd_sc_hd__a21o_1 _40001_ (.A1(_17416_),
    .A2(_17417_),
    .B1(_17418_),
    .X(_17419_));
 sky130_fd_sc_hd__nand3_4 _40002_ (.A(_17416_),
    .B(_17418_),
    .C(_17417_),
    .Y(_17420_));
 sky130_fd_sc_hd__o21ai_2 _40003_ (.A1(_17277_),
    .A2(_17278_),
    .B1(_17281_),
    .Y(_17421_));
 sky130_fd_sc_hd__a21oi_4 _40004_ (.A1(_17419_),
    .A2(_17420_),
    .B1(_17421_),
    .Y(_17422_));
 sky130_fd_sc_hd__and3_1 _40005_ (.A(_17419_),
    .B(_17421_),
    .C(_17420_),
    .X(_17423_));
 sky130_fd_sc_hd__nand2_1 _40006_ (.A(_19833_),
    .B(_20095_),
    .Y(_17424_));
 sky130_fd_sc_hd__and4_2 _40007_ (.A(_12604_),
    .B(_13837_),
    .C(_19830_),
    .D(_12304_),
    .X(_17425_));
 sky130_fd_sc_hd__o22a_1 _40008_ (.A1(_12303_),
    .A2(_11275_),
    .B1(_16102_),
    .B2(_08888_),
    .X(_17426_));
 sky130_fd_sc_hd__or3_4 _40009_ (.A(_17424_),
    .B(_17425_),
    .C(_17426_),
    .X(_17427_));
 sky130_fd_sc_hd__o21ai_2 _40010_ (.A1(_17425_),
    .A2(_17426_),
    .B1(_17424_),
    .Y(_17428_));
 sky130_fd_sc_hd__o21bai_2 _40011_ (.A1(_17245_),
    .A2(_17247_),
    .B1_N(_17246_),
    .Y(_17429_));
 sky130_fd_sc_hd__nand3_4 _40012_ (.A(_17427_),
    .B(_17428_),
    .C(_17429_),
    .Y(_17430_));
 sky130_fd_sc_hd__a21o_1 _40013_ (.A1(_17427_),
    .A2(_17428_),
    .B1(_17429_),
    .X(_17431_));
 sky130_fd_sc_hd__nand2_1 _40014_ (.A(_19845_),
    .B(_20084_),
    .Y(_17432_));
 sky130_fd_sc_hd__nor2_1 _40015_ (.A(_12307_),
    .B(_11941_),
    .Y(_17433_));
 sky130_fd_sc_hd__o22a_1 _40016_ (.A1(_16094_),
    .A2(_10781_),
    .B1(_16095_),
    .B2(_12307_),
    .X(_17434_));
 sky130_fd_sc_hd__a21o_1 _40017_ (.A1(_16093_),
    .A2(_17433_),
    .B1(_17434_),
    .X(_17435_));
 sky130_fd_sc_hd__nor2_4 _40018_ (.A(_17432_),
    .B(_17435_),
    .Y(_17436_));
 sky130_fd_sc_hd__and2_1 _40019_ (.A(_17435_),
    .B(_17432_),
    .X(_17437_));
 sky130_fd_sc_hd__o2bb2ai_4 _40020_ (.A1_N(_17430_),
    .A2_N(_17431_),
    .B1(_17436_),
    .B2(_17437_),
    .Y(_17438_));
 sky130_fd_sc_hd__nor2_2 _40021_ (.A(_17436_),
    .B(_17437_),
    .Y(_17439_));
 sky130_fd_sc_hd__nand3_4 _40022_ (.A(_17431_),
    .B(_17439_),
    .C(_17430_),
    .Y(_17440_));
 sky130_fd_sc_hd__a21o_1 _40023_ (.A1(_17269_),
    .A2(_17254_),
    .B1(_17253_),
    .X(_17441_));
 sky130_fd_sc_hd__a21oi_2 _40024_ (.A1(_17438_),
    .A2(_17440_),
    .B1(_17441_),
    .Y(_17442_));
 sky130_fd_sc_hd__nand2_1 _40025_ (.A(_17267_),
    .B(_17261_),
    .Y(_17443_));
 sky130_fd_sc_hd__o2111a_1 _40026_ (.A1(_17265_),
    .A2(_17266_),
    .B1(_17440_),
    .C1(_17443_),
    .D1(_17438_),
    .X(_17444_));
 sky130_fd_sc_hd__o22ai_4 _40027_ (.A1(_17422_),
    .A2(_17423_),
    .B1(_17442_),
    .B2(_17444_),
    .Y(_17445_));
 sky130_fd_sc_hd__a21o_1 _40028_ (.A1(_17438_),
    .A2(_17440_),
    .B1(_17441_),
    .X(_17446_));
 sky130_fd_sc_hd__nor2_2 _40029_ (.A(_17422_),
    .B(_17423_),
    .Y(_17447_));
 sky130_fd_sc_hd__nand3_4 _40030_ (.A(_17441_),
    .B(_17438_),
    .C(_17440_),
    .Y(_17448_));
 sky130_fd_sc_hd__nand3_4 _40031_ (.A(_17446_),
    .B(_17447_),
    .C(_17448_),
    .Y(_17449_));
 sky130_fd_sc_hd__nand2_1 _40032_ (.A(_17275_),
    .B(_17293_),
    .Y(_17450_));
 sky130_fd_sc_hd__nand2_2 _40033_ (.A(_17450_),
    .B(_17271_),
    .Y(_17451_));
 sky130_fd_sc_hd__a21oi_2 _40034_ (.A1(_17445_),
    .A2(_17449_),
    .B1(_17451_),
    .Y(_17452_));
 sky130_fd_sc_hd__and3_1 _40035_ (.A(_17262_),
    .B(_17264_),
    .C(_17270_),
    .X(_17453_));
 sky130_fd_sc_hd__a32oi_1 _40036_ (.A1(_17272_),
    .A2(_17273_),
    .A3(_17274_),
    .B1(_17292_),
    .B2(_17291_),
    .Y(_17454_));
 sky130_fd_sc_hd__o211a_1 _40037_ (.A1(_17453_),
    .A2(_17454_),
    .B1(_17449_),
    .C1(_17445_),
    .X(_17455_));
 sky130_fd_sc_hd__o22ai_4 _40038_ (.A1(_17409_),
    .A2(_17410_),
    .B1(_17452_),
    .B2(_17455_),
    .Y(_17456_));
 sky130_fd_sc_hd__a21o_1 _40039_ (.A1(_17445_),
    .A2(_17449_),
    .B1(_17451_),
    .X(_17457_));
 sky130_fd_sc_hd__nand3_2 _40040_ (.A(_17451_),
    .B(_17445_),
    .C(_17449_),
    .Y(_17458_));
 sky130_fd_sc_hd__nor2_2 _40041_ (.A(_17410_),
    .B(_17409_),
    .Y(_17459_));
 sky130_fd_sc_hd__nand3_4 _40042_ (.A(_17457_),
    .B(_17458_),
    .C(_17459_),
    .Y(_17460_));
 sky130_fd_sc_hd__o21ai_4 _40043_ (.A1(_17311_),
    .A2(_17297_),
    .B1(_17304_),
    .Y(_17461_));
 sky130_fd_sc_hd__a21oi_4 _40044_ (.A1(_17456_),
    .A2(_17460_),
    .B1(_17461_),
    .Y(_17462_));
 sky130_fd_sc_hd__a21oi_1 _40045_ (.A1(_17300_),
    .A2(_17301_),
    .B1(_17311_),
    .Y(_17463_));
 sky130_fd_sc_hd__o211a_2 _40046_ (.A1(_17298_),
    .A2(_17463_),
    .B1(_17460_),
    .C1(_17456_),
    .X(_17464_));
 sky130_fd_sc_hd__o22ai_4 _40047_ (.A1(_17394_),
    .A2(_17395_),
    .B1(_17462_),
    .B2(_17464_),
    .Y(_17465_));
 sky130_fd_sc_hd__a21o_1 _40048_ (.A1(_17456_),
    .A2(_17460_),
    .B1(_17461_),
    .X(_17466_));
 sky130_fd_sc_hd__nor2_4 _40049_ (.A(_17394_),
    .B(_17395_),
    .Y(_17467_));
 sky130_fd_sc_hd__nand3_2 _40050_ (.A(_17456_),
    .B(_17461_),
    .C(_17460_),
    .Y(_17468_));
 sky130_fd_sc_hd__nand3_2 _40051_ (.A(_17466_),
    .B(_17467_),
    .C(_17468_),
    .Y(_17469_));
 sky130_vsdinv _40052_ (.A(_17305_),
    .Y(_17470_));
 sky130_fd_sc_hd__nand2_1 _40053_ (.A(_17299_),
    .B(_17306_),
    .Y(_17471_));
 sky130_fd_sc_hd__o2bb2ai_2 _40054_ (.A1_N(_17331_),
    .A2_N(_17313_),
    .B1(_17470_),
    .B2(_17471_),
    .Y(_17472_));
 sky130_fd_sc_hd__nand3_4 _40055_ (.A(_17465_),
    .B(_17469_),
    .C(_17472_),
    .Y(_17473_));
 sky130_fd_sc_hd__o21ai_2 _40056_ (.A1(_17462_),
    .A2(_17464_),
    .B1(_17467_),
    .Y(_17474_));
 sky130_fd_sc_hd__a21boi_2 _40057_ (.A1(_17313_),
    .A2(_17331_),
    .B1_N(_17307_),
    .Y(_17475_));
 sky130_fd_sc_hd__nand3b_2 _40058_ (.A_N(_17467_),
    .B(_17466_),
    .C(_17468_),
    .Y(_17476_));
 sky130_fd_sc_hd__nand3_4 _40059_ (.A(_17474_),
    .B(_17475_),
    .C(_17476_),
    .Y(_17477_));
 sky130_fd_sc_hd__nor2_1 _40060_ (.A(_17323_),
    .B(_17322_),
    .Y(_17478_));
 sky130_fd_sc_hd__o21ai_2 _40061_ (.A1(_17325_),
    .A2(_17478_),
    .B1(_17324_),
    .Y(_17479_));
 sky130_fd_sc_hd__nor2_4 _40062_ (.A(_16783_),
    .B(_17479_),
    .Y(_17480_));
 sky130_fd_sc_hd__and2_2 _40063_ (.A(_17479_),
    .B(_16256_),
    .X(_17481_));
 sky130_fd_sc_hd__nor2_2 _40064_ (.A(_17480_),
    .B(_17481_),
    .Y(_17482_));
 sky130_fd_sc_hd__o21a_1 _40065_ (.A1(_16252_),
    .A2(_16255_),
    .B1(_17482_),
    .X(_17483_));
 sky130_fd_sc_hd__nor2_4 _40066_ (.A(_16787_),
    .B(_17482_),
    .Y(_17484_));
 sky130_fd_sc_hd__o2bb2ai_4 _40067_ (.A1_N(_17473_),
    .A2_N(_17477_),
    .B1(_17483_),
    .B2(_17484_),
    .Y(_17485_));
 sky130_fd_sc_hd__nor2_2 _40068_ (.A(_17484_),
    .B(_17483_),
    .Y(_17486_));
 sky130_fd_sc_hd__nand3_4 _40069_ (.A(_17486_),
    .B(_17477_),
    .C(_17473_),
    .Y(_17487_));
 sky130_fd_sc_hd__o21ai_4 _40070_ (.A1(_17344_),
    .A2(_17334_),
    .B1(_17351_),
    .Y(_17488_));
 sky130_fd_sc_hd__a21oi_4 _40071_ (.A1(_17485_),
    .A2(_17487_),
    .B1(_17488_),
    .Y(_17489_));
 sky130_fd_sc_hd__a21oi_1 _40072_ (.A1(_17348_),
    .A2(_17349_),
    .B1(_17344_),
    .Y(_17490_));
 sky130_fd_sc_hd__o211a_1 _40073_ (.A1(_17337_),
    .A2(_17490_),
    .B1(_17487_),
    .C1(_17485_),
    .X(_17491_));
 sky130_fd_sc_hd__nand2_1 _40074_ (.A(_17338_),
    .B(_16787_),
    .Y(_17492_));
 sky130_fd_sc_hd__nand2_1 _40075_ (.A(_17492_),
    .B(_17340_),
    .Y(_17493_));
 sky130_fd_sc_hd__nor2_1 _40076_ (.A(_14354_),
    .B(_17493_),
    .Y(_17494_));
 sky130_vsdinv _40077_ (.A(_17493_),
    .Y(_17495_));
 sky130_fd_sc_hd__nor2_1 _40078_ (.A(_16423_),
    .B(_17495_),
    .Y(_17496_));
 sky130_fd_sc_hd__nor2_2 _40079_ (.A(_17494_),
    .B(_17496_),
    .Y(_17497_));
 sky130_vsdinv _40080_ (.A(_17497_),
    .Y(_17498_));
 sky130_fd_sc_hd__o21ai_2 _40081_ (.A1(_17489_),
    .A2(_17491_),
    .B1(_17498_),
    .Y(_17499_));
 sky130_fd_sc_hd__a21boi_2 _40082_ (.A1(_17361_),
    .A2(_17367_),
    .B1_N(_17353_),
    .Y(_17500_));
 sky130_fd_sc_hd__a21o_1 _40083_ (.A1(_17485_),
    .A2(_17487_),
    .B1(_17488_),
    .X(_17501_));
 sky130_fd_sc_hd__nand3_4 _40084_ (.A(_17485_),
    .B(_17488_),
    .C(_17487_),
    .Y(_17502_));
 sky130_fd_sc_hd__nand3_2 _40085_ (.A(_17501_),
    .B(_17502_),
    .C(_17497_),
    .Y(_17503_));
 sky130_fd_sc_hd__nand3_4 _40086_ (.A(_17499_),
    .B(_17500_),
    .C(_17503_),
    .Y(_17504_));
 sky130_fd_sc_hd__o21ai_2 _40087_ (.A1(_17489_),
    .A2(_17491_),
    .B1(_17497_),
    .Y(_17505_));
 sky130_fd_sc_hd__nand3_2 _40088_ (.A(_17501_),
    .B(_17502_),
    .C(_17498_),
    .Y(_17506_));
 sky130_fd_sc_hd__nand2_1 _40089_ (.A(_17361_),
    .B(_17367_),
    .Y(_17507_));
 sky130_fd_sc_hd__nand2_1 _40090_ (.A(_17507_),
    .B(_17353_),
    .Y(_17508_));
 sky130_fd_sc_hd__nand3_4 _40091_ (.A(_17505_),
    .B(_17506_),
    .C(_17508_),
    .Y(_17509_));
 sky130_fd_sc_hd__a21o_2 _40092_ (.A1(_17504_),
    .A2(_17509_),
    .B1(_17366_),
    .X(_17510_));
 sky130_fd_sc_hd__nand3_4 _40093_ (.A(_17504_),
    .B(_17509_),
    .C(_17366_),
    .Y(_17511_));
 sky130_fd_sc_hd__nand2_1 _40094_ (.A(_17376_),
    .B(_17191_),
    .Y(_17512_));
 sky130_fd_sc_hd__nand2_4 _40095_ (.A(_17512_),
    .B(_17370_),
    .Y(_17513_));
 sky130_fd_sc_hd__a21oi_4 _40096_ (.A1(_17510_),
    .A2(_17511_),
    .B1(_17513_),
    .Y(_17514_));
 sky130_fd_sc_hd__and3_1 _40097_ (.A(_17510_),
    .B(_17511_),
    .C(_17513_),
    .X(_17515_));
 sky130_fd_sc_hd__nor2_4 _40098_ (.A(_17514_),
    .B(_17515_),
    .Y(_17516_));
 sky130_fd_sc_hd__nand3b_1 _40099_ (.A_N(_17386_),
    .B(_17384_),
    .C(_17516_),
    .Y(_17517_));
 sky130_vsdinv _40100_ (.A(_17384_),
    .Y(_17518_));
 sky130_fd_sc_hd__o21bai_1 _40101_ (.A1(_17518_),
    .A2(_17386_),
    .B1_N(_17516_),
    .Y(_17519_));
 sky130_fd_sc_hd__nand2_2 _40102_ (.A(_17517_),
    .B(_17519_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21o_1 _40103_ (.A1(_17466_),
    .A2(_17467_),
    .B1(_17464_),
    .X(_17520_));
 sky130_fd_sc_hd__nand2_2 _40104_ (.A(_17440_),
    .B(_17430_),
    .Y(_17521_));
 sky130_fd_sc_hd__nand2_1 _40105_ (.A(_16107_),
    .B(_20092_),
    .Y(_17522_));
 sky130_fd_sc_hd__or4_4 _40106_ (.A(_20099_),
    .B(_16448_),
    .C(_16102_),
    .D(_11557_),
    .X(_17523_));
 sky130_fd_sc_hd__a22o_1 _40107_ (.A1(_15907_),
    .A2(_20095_),
    .B1(_09880_),
    .B2(_15908_),
    .X(_17524_));
 sky130_fd_sc_hd__nand2_1 _40108_ (.A(_17523_),
    .B(_17524_),
    .Y(_17525_));
 sky130_fd_sc_hd__or2_2 _40109_ (.A(_17522_),
    .B(_17525_),
    .X(_17526_));
 sky130_fd_sc_hd__nand2_2 _40110_ (.A(_17525_),
    .B(_17522_),
    .Y(_17527_));
 sky130_fd_sc_hd__nand2_2 _40111_ (.A(_17526_),
    .B(_17527_),
    .Y(_17528_));
 sky130_vsdinv _40112_ (.A(_17425_),
    .Y(_17529_));
 sky130_fd_sc_hd__nand2_2 _40113_ (.A(_17427_),
    .B(_17529_),
    .Y(_17530_));
 sky130_vsdinv _40114_ (.A(_17530_),
    .Y(_17531_));
 sky130_fd_sc_hd__nand2_4 _40115_ (.A(_17528_),
    .B(_17531_),
    .Y(_17532_));
 sky130_fd_sc_hd__nand3_4 _40116_ (.A(_17526_),
    .B(_17530_),
    .C(_17527_),
    .Y(_17533_));
 sky130_fd_sc_hd__nand2_1 _40117_ (.A(_19845_),
    .B(_20080_),
    .Y(_17534_));
 sky130_fd_sc_hd__a22o_1 _40118_ (.A1(_15924_),
    .A2(_20087_),
    .B1(_15925_),
    .B2(_20083_),
    .X(_17535_));
 sky130_fd_sc_hd__o21ai_1 _40119_ (.A1(_16311_),
    .A2(_15867_),
    .B1(_17535_),
    .Y(_17536_));
 sky130_fd_sc_hd__or2_2 _40120_ (.A(_17534_),
    .B(_17536_),
    .X(_17537_));
 sky130_fd_sc_hd__nand2_1 _40121_ (.A(_17536_),
    .B(_17534_),
    .Y(_17538_));
 sky130_fd_sc_hd__nand2_2 _40122_ (.A(_17537_),
    .B(_17538_),
    .Y(_17539_));
 sky130_fd_sc_hd__nand3_2 _40123_ (.A(_17532_),
    .B(_17533_),
    .C(_17539_),
    .Y(_17540_));
 sky130_fd_sc_hd__nand2_1 _40124_ (.A(_17528_),
    .B(_17530_),
    .Y(_17541_));
 sky130_fd_sc_hd__nand3_2 _40125_ (.A(_17526_),
    .B(_17531_),
    .C(_17527_),
    .Y(_17542_));
 sky130_vsdinv _40126_ (.A(_17539_),
    .Y(_17543_));
 sky130_fd_sc_hd__nand3_2 _40127_ (.A(_17541_),
    .B(_17542_),
    .C(_17543_),
    .Y(_17544_));
 sky130_fd_sc_hd__nand3b_4 _40128_ (.A_N(_17521_),
    .B(_17540_),
    .C(_17544_),
    .Y(_17545_));
 sky130_fd_sc_hd__nand3_4 _40129_ (.A(_17532_),
    .B(_17533_),
    .C(_17543_),
    .Y(_17546_));
 sky130_fd_sc_hd__nand3_2 _40130_ (.A(_17541_),
    .B(_17542_),
    .C(_17539_),
    .Y(_17547_));
 sky130_fd_sc_hd__nand3_4 _40131_ (.A(_17546_),
    .B(_17547_),
    .C(_17521_),
    .Y(_17548_));
 sky130_fd_sc_hd__nand2_1 _40132_ (.A(_19852_),
    .B(_11604_),
    .Y(_17549_));
 sky130_fd_sc_hd__or3_4 _40133_ (.A(_17549_),
    .B(_16670_),
    .C(_10767_),
    .X(_17550_));
 sky130_fd_sc_hd__o21ai_2 _40134_ (.A1(_16670_),
    .A2(_16059_),
    .B1(_17549_),
    .Y(_17551_));
 sky130_fd_sc_hd__nor2_4 _40135_ (.A(_13024_),
    .B(net464),
    .Y(_17552_));
 sky130_fd_sc_hd__a21o_1 _40136_ (.A1(_17550_),
    .A2(_17551_),
    .B1(_17552_),
    .X(_17553_));
 sky130_fd_sc_hd__nand3_2 _40137_ (.A(_17550_),
    .B(_17552_),
    .C(_17551_),
    .Y(_17554_));
 sky130_fd_sc_hd__and2_1 _40138_ (.A(_17553_),
    .B(_17554_),
    .X(_17555_));
 sky130_fd_sc_hd__a21o_1 _40139_ (.A1(_16093_),
    .A2(_17433_),
    .B1(_17436_),
    .X(_17556_));
 sky130_fd_sc_hd__nor2_2 _40140_ (.A(_17555_),
    .B(_17556_),
    .Y(_17557_));
 sky130_fd_sc_hd__and2_1 _40141_ (.A(_17556_),
    .B(_17555_),
    .X(_17558_));
 sky130_fd_sc_hd__or3_4 _40142_ (.A(_17411_),
    .B(_15010_),
    .C(_16059_),
    .X(_17559_));
 sky130_fd_sc_hd__nand2_1 _40143_ (.A(_17416_),
    .B(_17559_),
    .Y(_17560_));
 sky130_fd_sc_hd__o21ai_2 _40144_ (.A1(_17557_),
    .A2(_17558_),
    .B1(_17560_),
    .Y(_17561_));
 sky130_vsdinv _40145_ (.A(_17560_),
    .Y(_17562_));
 sky130_fd_sc_hd__nand2_2 _40146_ (.A(_17556_),
    .B(_17555_),
    .Y(_17563_));
 sky130_fd_sc_hd__nand3b_2 _40147_ (.A_N(_17557_),
    .B(_17562_),
    .C(_17563_),
    .Y(_17564_));
 sky130_fd_sc_hd__nand2_4 _40148_ (.A(_17561_),
    .B(_17564_),
    .Y(_17565_));
 sky130_fd_sc_hd__a21o_1 _40149_ (.A1(_17545_),
    .A2(_17548_),
    .B1(_17565_),
    .X(_17566_));
 sky130_fd_sc_hd__nand3_4 _40150_ (.A(_17545_),
    .B(_17548_),
    .C(_17565_),
    .Y(_17567_));
 sky130_fd_sc_hd__nand2_2 _40151_ (.A(_17449_),
    .B(_17448_),
    .Y(_17568_));
 sky130_fd_sc_hd__a21o_1 _40152_ (.A1(_17566_),
    .A2(_17567_),
    .B1(_17568_),
    .X(_17569_));
 sky130_fd_sc_hd__nand3_4 _40153_ (.A(_17566_),
    .B(_17568_),
    .C(_17567_),
    .Y(_17570_));
 sky130_vsdinv _40154_ (.A(_19860_),
    .Y(_17571_));
 sky130_fd_sc_hd__or3_4 _40155_ (.A(_17221_),
    .B(_17571_),
    .C(_07822_),
    .X(_17572_));
 sky130_fd_sc_hd__nand2_1 _40156_ (.A(_17572_),
    .B(_17399_),
    .Y(_17573_));
 sky130_fd_sc_hd__or2_1 _40157_ (.A(_17573_),
    .B(_16884_),
    .X(_17574_));
 sky130_fd_sc_hd__nand2_1 _40158_ (.A(_16884_),
    .B(_17573_),
    .Y(_17575_));
 sky130_fd_sc_hd__and2_2 _40159_ (.A(_17574_),
    .B(_17575_),
    .X(_17576_));
 sky130_fd_sc_hd__a21bo_2 _40160_ (.A1(_17419_),
    .A2(_17421_),
    .B1_N(_17420_),
    .X(_17577_));
 sky130_fd_sc_hd__nand2_4 _40161_ (.A(_17576_),
    .B(_17577_),
    .Y(_17578_));
 sky130_vsdinv _40162_ (.A(_17572_),
    .Y(_17579_));
 sky130_fd_sc_hd__nor2_1 _40163_ (.A(_17579_),
    .B(_17401_),
    .Y(_17580_));
 sky130_vsdinv _40164_ (.A(_17580_),
    .Y(_17581_));
 sky130_fd_sc_hd__o21a_1 _40165_ (.A1(_17577_),
    .A2(_17576_),
    .B1(_17581_),
    .X(_17582_));
 sky130_fd_sc_hd__or2_1 _40166_ (.A(_17577_),
    .B(_17576_),
    .X(_17583_));
 sky130_fd_sc_hd__a21oi_2 _40167_ (.A1(_17583_),
    .A2(_17578_),
    .B1(_17581_),
    .Y(_17584_));
 sky130_fd_sc_hd__a21oi_4 _40168_ (.A1(_17578_),
    .A2(_17582_),
    .B1(_17584_),
    .Y(_17585_));
 sky130_fd_sc_hd__a21oi_2 _40169_ (.A1(_17569_),
    .A2(_17570_),
    .B1(_17585_),
    .Y(_17586_));
 sky130_fd_sc_hd__and3_1 _40170_ (.A(_17569_),
    .B(_17585_),
    .C(_17570_),
    .X(_17587_));
 sky130_fd_sc_hd__a21o_1 _40171_ (.A1(_17457_),
    .A2(_17459_),
    .B1(_17455_),
    .X(_17588_));
 sky130_fd_sc_hd__o21bai_4 _40172_ (.A1(_17586_),
    .A2(_17587_),
    .B1_N(_17588_),
    .Y(_17589_));
 sky130_fd_sc_hd__a21o_1 _40173_ (.A1(_17569_),
    .A2(_17570_),
    .B1(_17585_),
    .X(_17590_));
 sky130_fd_sc_hd__nand3_2 _40174_ (.A(_17569_),
    .B(_17585_),
    .C(_17570_),
    .Y(_17591_));
 sky130_fd_sc_hd__nand3_2 _40175_ (.A(_17590_),
    .B(_17591_),
    .C(_17588_),
    .Y(_17592_));
 sky130_fd_sc_hd__clkbuf_4 _40176_ (.A(_17592_),
    .X(_17593_));
 sky130_fd_sc_hd__buf_2 _40177_ (.A(_17393_),
    .X(_17594_));
 sky130_fd_sc_hd__nor2_1 _40178_ (.A(_17406_),
    .B(_17403_),
    .Y(_17595_));
 sky130_fd_sc_hd__nand2_1 _40179_ (.A(_17403_),
    .B(_17406_),
    .Y(_17596_));
 sky130_fd_sc_hd__o21ai_2 _40180_ (.A1(_17408_),
    .A2(_17595_),
    .B1(_17596_),
    .Y(_17597_));
 sky130_fd_sc_hd__or2_1 _40181_ (.A(_17323_),
    .B(_17597_),
    .X(_17598_));
 sky130_fd_sc_hd__nand2_2 _40182_ (.A(_17597_),
    .B(_17323_),
    .Y(_17599_));
 sky130_fd_sc_hd__nand2_2 _40183_ (.A(_17598_),
    .B(_17599_),
    .Y(_17600_));
 sky130_fd_sc_hd__nor2_1 _40184_ (.A(_17594_),
    .B(_17600_),
    .Y(_17601_));
 sky130_fd_sc_hd__nand2_1 _40185_ (.A(_17600_),
    .B(_17594_),
    .Y(_17602_));
 sky130_fd_sc_hd__and2b_1 _40186_ (.A_N(_17601_),
    .B(_17602_),
    .X(_17603_));
 sky130_fd_sc_hd__a21o_1 _40187_ (.A1(_17589_),
    .A2(_17593_),
    .B1(_17603_),
    .X(_17604_));
 sky130_fd_sc_hd__nand3_2 _40188_ (.A(_17589_),
    .B(_17593_),
    .C(_17603_),
    .Y(_17605_));
 sky130_fd_sc_hd__nand3b_4 _40189_ (.A_N(_17520_),
    .B(_17604_),
    .C(_17605_),
    .Y(_17606_));
 sky130_fd_sc_hd__or2b_4 _40190_ (.A(_17601_),
    .B_N(_17602_),
    .X(_17607_));
 sky130_fd_sc_hd__a21o_1 _40191_ (.A1(_17589_),
    .A2(_17592_),
    .B1(_17607_),
    .X(_17608_));
 sky130_fd_sc_hd__nand3_4 _40192_ (.A(_17589_),
    .B(_17593_),
    .C(_17607_),
    .Y(_17609_));
 sky130_fd_sc_hd__nand3_2 _40193_ (.A(_17608_),
    .B(_17609_),
    .C(_17520_),
    .Y(_17610_));
 sky130_fd_sc_hd__nand2_1 _40194_ (.A(_17606_),
    .B(_17610_),
    .Y(_17611_));
 sky130_fd_sc_hd__a21bo_1 _40195_ (.A1(_17388_),
    .A2(_17393_),
    .B1_N(_17390_),
    .X(_17612_));
 sky130_fd_sc_hd__clkbuf_4 _40196_ (.A(_16783_),
    .X(_17613_));
 sky130_fd_sc_hd__and2_2 _40197_ (.A(_17612_),
    .B(_17613_),
    .X(_17614_));
 sky130_vsdinv _40198_ (.A(_17614_),
    .Y(_17615_));
 sky130_fd_sc_hd__nor2_4 _40199_ (.A(_17613_),
    .B(_17612_),
    .Y(_17616_));
 sky130_fd_sc_hd__nor2_8 _40200_ (.A(_16982_),
    .B(_17616_),
    .Y(_17617_));
 sky130_fd_sc_hd__nor2_1 _40201_ (.A(_17616_),
    .B(_17614_),
    .Y(_17618_));
 sky130_fd_sc_hd__nor2_2 _40202_ (.A(_16975_),
    .B(_17618_),
    .Y(_17619_));
 sky130_fd_sc_hd__a21oi_4 _40203_ (.A1(_17615_),
    .A2(_17617_),
    .B1(_17619_),
    .Y(_17620_));
 sky130_fd_sc_hd__nand2_1 _40204_ (.A(_17611_),
    .B(_17620_),
    .Y(_17621_));
 sky130_fd_sc_hd__nand2_2 _40205_ (.A(_17487_),
    .B(_17473_),
    .Y(_17622_));
 sky130_vsdinv _40206_ (.A(_17622_),
    .Y(_17623_));
 sky130_fd_sc_hd__buf_4 _40207_ (.A(_17610_),
    .X(_17624_));
 sky130_fd_sc_hd__a21o_1 _40208_ (.A1(_17615_),
    .A2(_17617_),
    .B1(_17619_),
    .X(_17625_));
 sky130_fd_sc_hd__nand3_2 _40209_ (.A(_17606_),
    .B(_17624_),
    .C(_17625_),
    .Y(_17626_));
 sky130_fd_sc_hd__nand3_4 _40210_ (.A(_17621_),
    .B(_17623_),
    .C(_17626_),
    .Y(_17627_));
 sky130_fd_sc_hd__nand2_1 _40211_ (.A(_17611_),
    .B(_17625_),
    .Y(_17628_));
 sky130_fd_sc_hd__nand3_2 _40212_ (.A(_17606_),
    .B(_17624_),
    .C(_17620_),
    .Y(_17629_));
 sky130_fd_sc_hd__nand3_4 _40213_ (.A(_17628_),
    .B(_17622_),
    .C(_17629_),
    .Y(_17630_));
 sky130_fd_sc_hd__nor2_4 _40214_ (.A(_16992_),
    .B(_17480_),
    .Y(_17631_));
 sky130_fd_sc_hd__nor2_8 _40215_ (.A(_17481_),
    .B(_17631_),
    .Y(_17632_));
 sky130_fd_sc_hd__buf_4 _40216_ (.A(_16426_),
    .X(_17633_));
 sky130_fd_sc_hd__and2_1 _40217_ (.A(_17632_),
    .B(_17633_),
    .X(_17634_));
 sky130_fd_sc_hd__nor2_1 _40218_ (.A(_17633_),
    .B(_17632_),
    .Y(_17635_));
 sky130_fd_sc_hd__o2bb2ai_2 _40219_ (.A1_N(_17627_),
    .A2_N(_17630_),
    .B1(_17634_),
    .B2(_17635_),
    .Y(_17636_));
 sky130_fd_sc_hd__nand2_1 _40220_ (.A(_17501_),
    .B(_17498_),
    .Y(_17637_));
 sky130_fd_sc_hd__nand2_2 _40221_ (.A(_17637_),
    .B(_17502_),
    .Y(_17638_));
 sky130_vsdinv _40222_ (.A(_17638_),
    .Y(_17639_));
 sky130_fd_sc_hd__nor2_8 _40223_ (.A(_14355_),
    .B(_17632_),
    .Y(_17640_));
 sky130_fd_sc_hd__nand2_1 _40224_ (.A(_17632_),
    .B(net413),
    .Y(_17641_));
 sky130_vsdinv _40225_ (.A(_17641_),
    .Y(_17642_));
 sky130_fd_sc_hd__nor2_4 _40226_ (.A(_17640_),
    .B(_17642_),
    .Y(_17643_));
 sky130_fd_sc_hd__nand3b_4 _40227_ (.A_N(_17643_),
    .B(_17630_),
    .C(_17627_),
    .Y(_17644_));
 sky130_fd_sc_hd__nand3_2 _40228_ (.A(_17636_),
    .B(_17639_),
    .C(_17644_),
    .Y(_17645_));
 sky130_fd_sc_hd__o2bb2ai_2 _40229_ (.A1_N(_17627_),
    .A2_N(_17630_),
    .B1(_17640_),
    .B2(_17642_),
    .Y(_17646_));
 sky130_fd_sc_hd__nand3_2 _40230_ (.A(_17630_),
    .B(_17627_),
    .C(_17643_),
    .Y(_17647_));
 sky130_fd_sc_hd__nand3_4 _40231_ (.A(_17646_),
    .B(_17638_),
    .C(_17647_),
    .Y(_17648_));
 sky130_fd_sc_hd__nor2_2 _40232_ (.A(_16818_),
    .B(_17495_),
    .Y(_17649_));
 sky130_fd_sc_hd__a21oi_1 _40233_ (.A1(_17645_),
    .A2(_17648_),
    .B1(_17649_),
    .Y(_17650_));
 sky130_fd_sc_hd__and3_1 _40234_ (.A(_17648_),
    .B(_17645_),
    .C(_17649_),
    .X(_17651_));
 sky130_fd_sc_hd__nand2_2 _40235_ (.A(_17511_),
    .B(_17509_),
    .Y(_17652_));
 sky130_fd_sc_hd__o21bai_1 _40236_ (.A1(_17650_),
    .A2(_17651_),
    .B1_N(_17652_),
    .Y(_17653_));
 sky130_fd_sc_hd__a21o_1 _40237_ (.A1(_17645_),
    .A2(_17648_),
    .B1(_17649_),
    .X(_17654_));
 sky130_vsdinv _40238_ (.A(_17649_),
    .Y(_17655_));
 sky130_fd_sc_hd__a31oi_4 _40239_ (.A1(_17636_),
    .A2(_17639_),
    .A3(_17644_),
    .B1(_17655_),
    .Y(_17656_));
 sky130_fd_sc_hd__nand2_1 _40240_ (.A(_17656_),
    .B(_17648_),
    .Y(_17657_));
 sky130_fd_sc_hd__nand3_4 _40241_ (.A(_17654_),
    .B(_17652_),
    .C(_17657_),
    .Y(_17658_));
 sky130_fd_sc_hd__and2_1 _40242_ (.A(_17653_),
    .B(_17658_),
    .X(_17659_));
 sky130_fd_sc_hd__nand3_2 _40243_ (.A(_17211_),
    .B(_17516_),
    .C(_17385_),
    .Y(_17660_));
 sky130_fd_sc_hd__nand3_4 _40244_ (.A(_17510_),
    .B(_17511_),
    .C(_17513_),
    .Y(_17661_));
 sky130_fd_sc_hd__o21ai_2 _40245_ (.A1(_17384_),
    .A2(_17514_),
    .B1(_17661_),
    .Y(_17662_));
 sky130_fd_sc_hd__a31oi_4 _40246_ (.A1(_17516_),
    .A2(_17385_),
    .A3(_17214_),
    .B1(_17662_),
    .Y(_17663_));
 sky130_fd_sc_hd__o21ai_4 _40247_ (.A1(_17660_),
    .A2(_17028_),
    .B1(_17663_),
    .Y(_17664_));
 sky130_fd_sc_hd__o2111ai_4 _40248_ (.A1(_17208_),
    .A2(_17210_),
    .B1(_17022_),
    .C1(_17205_),
    .D1(_17016_),
    .Y(_17665_));
 sky130_fd_sc_hd__nand2_1 _40249_ (.A(_17382_),
    .B(_17380_),
    .Y(_17666_));
 sky130_fd_sc_hd__a21oi_1 _40250_ (.A1(_17504_),
    .A2(_17509_),
    .B1(_17366_),
    .Y(_17667_));
 sky130_fd_sc_hd__and3_1 _40251_ (.A(_17504_),
    .B(_17509_),
    .C(_17366_),
    .X(_17668_));
 sky130_fd_sc_hd__o21bai_2 _40252_ (.A1(_17667_),
    .A2(_17668_),
    .B1_N(_17513_),
    .Y(_17669_));
 sky130_fd_sc_hd__o2111ai_4 _40253_ (.A1(_17378_),
    .A2(_17666_),
    .B1(_17661_),
    .C1(_17381_),
    .D1(_17669_),
    .Y(_17670_));
 sky130_fd_sc_hd__nor2_1 _40254_ (.A(_17665_),
    .B(_17670_),
    .Y(_17671_));
 sky130_fd_sc_hd__nand2_1 _40255_ (.A(_17671_),
    .B(_17031_),
    .Y(_17672_));
 sky130_fd_sc_hd__a21oi_4 _40256_ (.A1(_16238_),
    .A2(_16241_),
    .B1(_17672_),
    .Y(_17673_));
 sky130_fd_sc_hd__or2_1 _40257_ (.A(_17664_),
    .B(_17673_),
    .X(_17674_));
 sky130_fd_sc_hd__or2_1 _40258_ (.A(_17659_),
    .B(_17674_),
    .X(_17675_));
 sky130_fd_sc_hd__nand2_1 _40259_ (.A(_17674_),
    .B(_17659_),
    .Y(_17676_));
 sky130_fd_sc_hd__and2_2 _40260_ (.A(_17675_),
    .B(_17676_),
    .X(_02675_));
 sky130_vsdinv _40261_ (.A(_17640_),
    .Y(_17677_));
 sky130_fd_sc_hd__nand2_2 _40262_ (.A(_17606_),
    .B(_17620_),
    .Y(_17678_));
 sky130_fd_sc_hd__nand2_1 _40263_ (.A(_17678_),
    .B(_17624_),
    .Y(_17679_));
 sky130_fd_sc_hd__a21boi_4 _40264_ (.A1(_17589_),
    .A2(_17607_),
    .B1_N(_17593_),
    .Y(_17680_));
 sky130_fd_sc_hd__a21boi_4 _40265_ (.A1(_17532_),
    .A2(_17543_),
    .B1_N(_17533_),
    .Y(_17681_));
 sky130_fd_sc_hd__o21a_2 _40266_ (.A1(_17522_),
    .A2(_17525_),
    .B1(_17523_),
    .X(_17682_));
 sky130_vsdinv _40267_ (.A(_17682_),
    .Y(_17683_));
 sky130_fd_sc_hd__nand2_2 _40268_ (.A(_19834_),
    .B(_20089_),
    .Y(_17684_));
 sky130_fd_sc_hd__or4_4 _40269_ (.A(_20095_),
    .B(_16448_),
    .C(_15916_),
    .D(_11941_),
    .X(_17685_));
 sky130_fd_sc_hd__a22o_1 _40270_ (.A1(_19831_),
    .A2(_20092_),
    .B1(_11563_),
    .B2(_15908_),
    .X(_17686_));
 sky130_fd_sc_hd__nand2_2 _40271_ (.A(_17685_),
    .B(_17686_),
    .Y(_17687_));
 sky130_fd_sc_hd__or2_4 _40272_ (.A(_17684_),
    .B(_17687_),
    .X(_17688_));
 sky130_fd_sc_hd__nand2_4 _40273_ (.A(_17687_),
    .B(_17684_),
    .Y(_17689_));
 sky130_fd_sc_hd__nand3_4 _40274_ (.A(_17683_),
    .B(_17688_),
    .C(_17689_),
    .Y(_17690_));
 sky130_fd_sc_hd__nand2_2 _40275_ (.A(_17688_),
    .B(_17689_),
    .Y(_17691_));
 sky130_fd_sc_hd__nand2_4 _40276_ (.A(_17691_),
    .B(_17682_),
    .Y(_17692_));
 sky130_fd_sc_hd__nand2_1 _40277_ (.A(_15897_),
    .B(_20075_),
    .Y(_17693_));
 sky130_fd_sc_hd__a22o_1 _40278_ (.A1(_19836_),
    .A2(_11165_),
    .B1(_15925_),
    .B2(_20079_),
    .X(_17694_));
 sky130_fd_sc_hd__o21ai_1 _40279_ (.A1(_10988_),
    .A2(_16056_),
    .B1(_17694_),
    .Y(_17695_));
 sky130_fd_sc_hd__or2_2 _40280_ (.A(_17693_),
    .B(_17695_),
    .X(_17696_));
 sky130_fd_sc_hd__nand2_1 _40281_ (.A(_17695_),
    .B(_17693_),
    .Y(_17697_));
 sky130_fd_sc_hd__nand2_4 _40282_ (.A(_17696_),
    .B(_17697_),
    .Y(_17698_));
 sky130_fd_sc_hd__nand3_2 _40283_ (.A(_17690_),
    .B(_17692_),
    .C(_17698_),
    .Y(_17699_));
 sky130_fd_sc_hd__nand2_2 _40284_ (.A(_17691_),
    .B(_17683_),
    .Y(_17700_));
 sky130_fd_sc_hd__nand3_4 _40285_ (.A(_17688_),
    .B(_17682_),
    .C(_17689_),
    .Y(_17701_));
 sky130_vsdinv _40286_ (.A(_17698_),
    .Y(_17702_));
 sky130_fd_sc_hd__nand3_2 _40287_ (.A(_17700_),
    .B(_17701_),
    .C(_17702_),
    .Y(_17703_));
 sky130_fd_sc_hd__nand3_4 _40288_ (.A(_17681_),
    .B(_17699_),
    .C(_17703_),
    .Y(_17704_));
 sky130_fd_sc_hd__nand2_2 _40289_ (.A(_17546_),
    .B(_17533_),
    .Y(_17705_));
 sky130_fd_sc_hd__nand3_4 _40290_ (.A(_17690_),
    .B(_17692_),
    .C(_17702_),
    .Y(_17706_));
 sky130_fd_sc_hd__nand3_4 _40291_ (.A(_17700_),
    .B(_17701_),
    .C(_17698_),
    .Y(_17707_));
 sky130_fd_sc_hd__nand3_4 _40292_ (.A(_17705_),
    .B(_17706_),
    .C(_17707_),
    .Y(_17708_));
 sky130_vsdinv _40293_ (.A(_17552_),
    .Y(_17709_));
 sky130_fd_sc_hd__nand2_8 _40294_ (.A(net503),
    .B(_10384_),
    .Y(_17710_));
 sky130_fd_sc_hd__or3_4 _40295_ (.A(_17710_),
    .B(_16670_),
    .C(_11176_),
    .X(_17711_));
 sky130_fd_sc_hd__o21ai_2 _40296_ (.A1(_16670_),
    .A2(_16147_),
    .B1(_17710_),
    .Y(_17712_));
 sky130_fd_sc_hd__nand2_1 _40297_ (.A(_17711_),
    .B(_17712_),
    .Y(_17713_));
 sky130_fd_sc_hd__or2_1 _40298_ (.A(_17709_),
    .B(_17713_),
    .X(_17714_));
 sky130_fd_sc_hd__nand2_1 _40299_ (.A(_17713_),
    .B(_17709_),
    .Y(_17715_));
 sky130_fd_sc_hd__and2_1 _40300_ (.A(_17714_),
    .B(_17715_),
    .X(_17716_));
 sky130_fd_sc_hd__o21ai_4 _40301_ (.A1(_16327_),
    .A2(_15867_),
    .B1(_17537_),
    .Y(_17717_));
 sky130_fd_sc_hd__nand2_4 _40302_ (.A(_17716_),
    .B(_17717_),
    .Y(_17718_));
 sky130_fd_sc_hd__a21o_2 _40303_ (.A1(_17714_),
    .A2(_17715_),
    .B1(_17717_),
    .X(_17719_));
 sky130_fd_sc_hd__nand2_4 _40304_ (.A(_17554_),
    .B(_17550_),
    .Y(_17720_));
 sky130_vsdinv _40305_ (.A(_17720_),
    .Y(_17721_));
 sky130_fd_sc_hd__a21oi_4 _40306_ (.A1(_17718_),
    .A2(_17719_),
    .B1(_17721_),
    .Y(_17722_));
 sky130_fd_sc_hd__nand2_2 _40307_ (.A(_17718_),
    .B(_17719_),
    .Y(_17723_));
 sky130_fd_sc_hd__nor2_4 _40308_ (.A(_17720_),
    .B(_17723_),
    .Y(_17724_));
 sky130_fd_sc_hd__o2bb2ai_2 _40309_ (.A1_N(_17704_),
    .A2_N(_17708_),
    .B1(_17722_),
    .B2(_17724_),
    .Y(_17725_));
 sky130_fd_sc_hd__a21boi_2 _40310_ (.A1(_17545_),
    .A2(_17565_),
    .B1_N(_17548_),
    .Y(_17726_));
 sky130_fd_sc_hd__a21oi_4 _40311_ (.A1(_17718_),
    .A2(_17719_),
    .B1(_17720_),
    .Y(_17727_));
 sky130_fd_sc_hd__nor2_4 _40312_ (.A(_17721_),
    .B(_17723_),
    .Y(_17728_));
 sky130_fd_sc_hd__o211ai_4 _40313_ (.A1(_17727_),
    .A2(_17728_),
    .B1(_17704_),
    .C1(_17708_),
    .Y(_17729_));
 sky130_fd_sc_hd__nand3_4 _40314_ (.A(_17725_),
    .B(_17726_),
    .C(_17729_),
    .Y(_17730_));
 sky130_fd_sc_hd__o2bb2ai_2 _40315_ (.A1_N(_17704_),
    .A2_N(_17708_),
    .B1(_17728_),
    .B2(_17727_),
    .Y(_17731_));
 sky130_fd_sc_hd__nand2_1 _40316_ (.A(_17567_),
    .B(_17548_),
    .Y(_17732_));
 sky130_fd_sc_hd__o211ai_4 _40317_ (.A1(_17722_),
    .A2(_17724_),
    .B1(_17704_),
    .C1(_17708_),
    .Y(_17733_));
 sky130_fd_sc_hd__nand3_4 _40318_ (.A(_17731_),
    .B(_17732_),
    .C(_17733_),
    .Y(_17734_));
 sky130_fd_sc_hd__nor2_8 _40319_ (.A(_17572_),
    .B(_16885_),
    .Y(_17735_));
 sky130_vsdinv _40320_ (.A(_17399_),
    .Y(_17736_));
 sky130_fd_sc_hd__nand2_2 _40321_ (.A(_16885_),
    .B(_17736_),
    .Y(_17737_));
 sky130_vsdinv _40322_ (.A(_17737_),
    .Y(_17738_));
 sky130_fd_sc_hd__nor2_8 _40323_ (.A(_17735_),
    .B(_17738_),
    .Y(_17739_));
 sky130_fd_sc_hd__a211o_1 _40324_ (.A1(_17559_),
    .A2(_17416_),
    .B1(_17557_),
    .C1(_17558_),
    .X(_17740_));
 sky130_fd_sc_hd__nand2_4 _40325_ (.A(_17740_),
    .B(_17563_),
    .Y(_17741_));
 sky130_fd_sc_hd__xor2_4 _40326_ (.A(_17739_),
    .B(_17741_),
    .X(_17742_));
 sky130_fd_sc_hd__a21o_1 _40327_ (.A1(_17730_),
    .A2(_17734_),
    .B1(_17742_),
    .X(_17743_));
 sky130_fd_sc_hd__a21o_1 _40328_ (.A1(_17583_),
    .A2(_17578_),
    .B1(_17581_),
    .X(_17744_));
 sky130_fd_sc_hd__nand2_2 _40329_ (.A(_17582_),
    .B(_17578_),
    .Y(_17745_));
 sky130_fd_sc_hd__nand2_1 _40330_ (.A(_17744_),
    .B(_17745_),
    .Y(_17746_));
 sky130_fd_sc_hd__a21oi_2 _40331_ (.A1(_17566_),
    .A2(_17567_),
    .B1(_17568_),
    .Y(_17747_));
 sky130_fd_sc_hd__o21ai_2 _40332_ (.A1(_17746_),
    .A2(_17747_),
    .B1(_17570_),
    .Y(_17748_));
 sky130_fd_sc_hd__nand3_4 _40333_ (.A(_17734_),
    .B(_17730_),
    .C(_17742_),
    .Y(_17749_));
 sky130_fd_sc_hd__nand3_4 _40334_ (.A(_17743_),
    .B(_17748_),
    .C(_17749_),
    .Y(_17750_));
 sky130_fd_sc_hd__a21oi_2 _40335_ (.A1(_17734_),
    .A2(_17730_),
    .B1(_17742_),
    .Y(_17751_));
 sky130_vsdinv _40336_ (.A(_17739_),
    .Y(_17752_));
 sky130_fd_sc_hd__nor2_1 _40337_ (.A(_17752_),
    .B(_17741_),
    .Y(_17753_));
 sky130_vsdinv _40338_ (.A(_17741_),
    .Y(_17754_));
 sky130_fd_sc_hd__nor2_1 _40339_ (.A(_17739_),
    .B(_17754_),
    .Y(_17755_));
 sky130_fd_sc_hd__o211a_1 _40340_ (.A1(_17753_),
    .A2(_17755_),
    .B1(_17730_),
    .C1(_17734_),
    .X(_17756_));
 sky130_fd_sc_hd__o21a_1 _40341_ (.A1(_17746_),
    .A2(_17747_),
    .B1(_17570_),
    .X(_17757_));
 sky130_fd_sc_hd__o21ai_4 _40342_ (.A1(_17751_),
    .A2(_17756_),
    .B1(_17757_),
    .Y(_17758_));
 sky130_fd_sc_hd__clkbuf_4 _40343_ (.A(_17391_),
    .X(_17759_));
 sky130_fd_sc_hd__a21o_1 _40344_ (.A1(_17745_),
    .A2(_17578_),
    .B1(_17320_),
    .X(_17760_));
 sky130_fd_sc_hd__nand3_4 _40345_ (.A(_17745_),
    .B(_17320_),
    .C(_17578_),
    .Y(_17761_));
 sky130_fd_sc_hd__nand2_1 _40346_ (.A(_17760_),
    .B(_17761_),
    .Y(_17762_));
 sky130_vsdinv _40347_ (.A(_17762_),
    .Y(_17763_));
 sky130_fd_sc_hd__nor2_2 _40348_ (.A(_17759_),
    .B(_17763_),
    .Y(_17764_));
 sky130_fd_sc_hd__clkbuf_4 _40349_ (.A(_17393_),
    .X(_17765_));
 sky130_fd_sc_hd__nor2_2 _40350_ (.A(_17765_),
    .B(_17762_),
    .Y(_17766_));
 sky130_fd_sc_hd__o2bb2ai_4 _40351_ (.A1_N(_17750_),
    .A2_N(_17758_),
    .B1(_17764_),
    .B2(_17766_),
    .Y(_17767_));
 sky130_fd_sc_hd__nand2_1 _40352_ (.A(_17762_),
    .B(_17391_),
    .Y(_17768_));
 sky130_fd_sc_hd__nand3_4 _40353_ (.A(_17760_),
    .B(_17393_),
    .C(_17761_),
    .Y(_17769_));
 sky130_fd_sc_hd__nand2_2 _40354_ (.A(_17768_),
    .B(_17769_),
    .Y(_17770_));
 sky130_fd_sc_hd__nand3_4 _40355_ (.A(_17758_),
    .B(_17750_),
    .C(_17770_),
    .Y(_17771_));
 sky130_fd_sc_hd__nand3_4 _40356_ (.A(_17680_),
    .B(_17767_),
    .C(_17771_),
    .Y(_17772_));
 sky130_fd_sc_hd__a21oi_2 _40357_ (.A1(_17590_),
    .A2(_17591_),
    .B1(_17588_),
    .Y(_17773_));
 sky130_fd_sc_hd__o21ai_2 _40358_ (.A1(_17603_),
    .A2(_17773_),
    .B1(_17593_),
    .Y(_17774_));
 sky130_vsdinv _40359_ (.A(_17769_),
    .Y(_17775_));
 sky130_vsdinv _40360_ (.A(_17768_),
    .Y(_17776_));
 sky130_fd_sc_hd__o2bb2ai_1 _40361_ (.A1_N(_17750_),
    .A2_N(_17758_),
    .B1(_17775_),
    .B2(_17776_),
    .Y(_17777_));
 sky130_fd_sc_hd__and2_1 _40362_ (.A(_17768_),
    .B(_17769_),
    .X(_17778_));
 sky130_fd_sc_hd__nand3_2 _40363_ (.A(_17758_),
    .B(_17778_),
    .C(_17750_),
    .Y(_17779_));
 sky130_fd_sc_hd__nand3_4 _40364_ (.A(_17774_),
    .B(_17777_),
    .C(_17779_),
    .Y(_17780_));
 sky130_fd_sc_hd__o21ai_1 _40365_ (.A1(_17391_),
    .A2(_17600_),
    .B1(_17599_),
    .Y(_17781_));
 sky130_fd_sc_hd__nand2_2 _40366_ (.A(_17781_),
    .B(_17613_),
    .Y(_17782_));
 sky130_vsdinv _40367_ (.A(_17782_),
    .Y(_17783_));
 sky130_fd_sc_hd__o211ai_4 _40368_ (.A1(_17759_),
    .A2(_17600_),
    .B1(_16971_),
    .C1(_17599_),
    .Y(_17784_));
 sky130_fd_sc_hd__nand2_2 _40369_ (.A(_17784_),
    .B(_16592_),
    .Y(_17785_));
 sky130_fd_sc_hd__nand2_2 _40370_ (.A(_17782_),
    .B(_17784_),
    .Y(_17786_));
 sky130_fd_sc_hd__nand2_2 _40371_ (.A(_17786_),
    .B(_16992_),
    .Y(_17787_));
 sky130_fd_sc_hd__o21a_2 _40372_ (.A1(_17783_),
    .A2(_17785_),
    .B1(_17787_),
    .X(_17788_));
 sky130_fd_sc_hd__a21o_1 _40373_ (.A1(_17772_),
    .A2(_17780_),
    .B1(_17788_),
    .X(_17789_));
 sky130_fd_sc_hd__nand3_2 _40374_ (.A(_17772_),
    .B(_17780_),
    .C(_17788_),
    .Y(_17790_));
 sky130_fd_sc_hd__nand3_4 _40375_ (.A(_17679_),
    .B(_17789_),
    .C(_17790_),
    .Y(_17791_));
 sky130_fd_sc_hd__a21oi_4 _40376_ (.A1(_17608_),
    .A2(_17609_),
    .B1(_17520_),
    .Y(_17792_));
 sky130_fd_sc_hd__o21ai_4 _40377_ (.A1(_17785_),
    .A2(_17783_),
    .B1(_17787_),
    .Y(_17793_));
 sky130_fd_sc_hd__nand3_4 _40378_ (.A(_17772_),
    .B(_17780_),
    .C(_17793_),
    .Y(_17794_));
 sky130_fd_sc_hd__and2_1 _40379_ (.A(_17786_),
    .B(_16975_),
    .X(_17795_));
 sky130_fd_sc_hd__clkbuf_4 _40380_ (.A(_16787_),
    .X(_17796_));
 sky130_fd_sc_hd__nor2_2 _40381_ (.A(_17796_),
    .B(_17786_),
    .Y(_17797_));
 sky130_fd_sc_hd__o2bb2ai_4 _40382_ (.A1_N(_17780_),
    .A2_N(_17772_),
    .B1(_17795_),
    .B2(_17797_),
    .Y(_17798_));
 sky130_fd_sc_hd__o2111ai_4 _40383_ (.A1(_17625_),
    .A2(_17792_),
    .B1(_17624_),
    .C1(_17794_),
    .D1(_17798_),
    .Y(_17799_));
 sky130_fd_sc_hd__nor3_4 _40384_ (.A(_16423_),
    .B(_17614_),
    .C(_17617_),
    .Y(_17800_));
 sky130_fd_sc_hd__o21a_1 _40385_ (.A1(_17614_),
    .A2(_17617_),
    .B1(_16423_),
    .X(_17801_));
 sky130_fd_sc_hd__nor2_2 _40386_ (.A(_17800_),
    .B(_17801_),
    .Y(_17802_));
 sky130_vsdinv _40387_ (.A(_17802_),
    .Y(_17803_));
 sky130_fd_sc_hd__a21o_1 _40388_ (.A1(_17791_),
    .A2(_17799_),
    .B1(_17803_),
    .X(_17804_));
 sky130_fd_sc_hd__a21boi_4 _40389_ (.A1(_17627_),
    .A2(_17643_),
    .B1_N(_17630_),
    .Y(_17805_));
 sky130_fd_sc_hd__nand3_4 _40390_ (.A(_17791_),
    .B(_17803_),
    .C(_17799_),
    .Y(_17806_));
 sky130_fd_sc_hd__nand3_2 _40391_ (.A(_17804_),
    .B(_17805_),
    .C(_17806_),
    .Y(_17807_));
 sky130_fd_sc_hd__nand2_1 _40392_ (.A(_17627_),
    .B(_17643_),
    .Y(_17808_));
 sky130_fd_sc_hd__nand2_1 _40393_ (.A(_17808_),
    .B(_17630_),
    .Y(_17809_));
 sky130_fd_sc_hd__clkbuf_2 _40394_ (.A(_17801_),
    .X(_17810_));
 sky130_fd_sc_hd__o2bb2ai_1 _40395_ (.A1_N(_17799_),
    .A2_N(_17791_),
    .B1(_17810_),
    .B2(_17800_),
    .Y(_17811_));
 sky130_fd_sc_hd__a41oi_4 _40396_ (.A1(_17624_),
    .A2(_17798_),
    .A3(_17678_),
    .A4(_17794_),
    .B1(_17803_),
    .Y(_17812_));
 sky130_fd_sc_hd__nand2_1 _40397_ (.A(_17812_),
    .B(_17791_),
    .Y(_17813_));
 sky130_fd_sc_hd__nand3_2 _40398_ (.A(_17809_),
    .B(_17811_),
    .C(_17813_),
    .Y(_17814_));
 sky130_fd_sc_hd__nand2_1 _40399_ (.A(_17807_),
    .B(_17814_),
    .Y(_17815_));
 sky130_fd_sc_hd__nor2_1 _40400_ (.A(_17677_),
    .B(_17815_),
    .Y(_17816_));
 sky130_vsdinv _40401_ (.A(_17648_),
    .Y(_17817_));
 sky130_fd_sc_hd__o2bb2ai_1 _40402_ (.A1_N(_17677_),
    .A2_N(_17815_),
    .B1(_17656_),
    .B2(_17817_),
    .Y(_17818_));
 sky130_fd_sc_hd__or2_2 _40403_ (.A(_17816_),
    .B(_17818_),
    .X(_17819_));
 sky130_fd_sc_hd__nor2_1 _40404_ (.A(_17656_),
    .B(_17817_),
    .Y(_17820_));
 sky130_fd_sc_hd__nand2_1 _40405_ (.A(_17815_),
    .B(_17640_),
    .Y(_17821_));
 sky130_fd_sc_hd__nand3_1 _40406_ (.A(_17807_),
    .B(_17814_),
    .C(_17677_),
    .Y(_17822_));
 sky130_fd_sc_hd__nand3_2 _40407_ (.A(_17820_),
    .B(_17821_),
    .C(_17822_),
    .Y(_17823_));
 sky130_fd_sc_hd__nand2_2 _40408_ (.A(_17819_),
    .B(_17823_),
    .Y(_17824_));
 sky130_fd_sc_hd__nand2_2 _40409_ (.A(_17676_),
    .B(_17658_),
    .Y(_17825_));
 sky130_fd_sc_hd__xnor2_4 _40410_ (.A(_17824_),
    .B(_17825_),
    .Y(_02676_));
 sky130_fd_sc_hd__o2111a_1 _40411_ (.A1(_17816_),
    .A2(_17818_),
    .B1(_17658_),
    .C1(_17823_),
    .D1(_17653_),
    .X(_17826_));
 sky130_fd_sc_hd__nand2_2 _40412_ (.A(_17674_),
    .B(_17826_),
    .Y(_17827_));
 sky130_vsdinv _40413_ (.A(_17823_),
    .Y(_17828_));
 sky130_fd_sc_hd__a21oi_4 _40414_ (.A1(_17819_),
    .A2(_17658_),
    .B1(_17828_),
    .Y(_17829_));
 sky130_vsdinv _40415_ (.A(_17829_),
    .Y(_17830_));
 sky130_fd_sc_hd__a22oi_4 _40416_ (.A1(_17678_),
    .A2(_17624_),
    .B1(_17798_),
    .B2(_17794_),
    .Y(_17831_));
 sky130_fd_sc_hd__a21o_1 _40417_ (.A1(_17741_),
    .A2(_17737_),
    .B1(_17735_),
    .X(_17832_));
 sky130_fd_sc_hd__buf_2 _40418_ (.A(_17319_),
    .X(_17833_));
 sky130_fd_sc_hd__nand2_2 _40419_ (.A(_17832_),
    .B(_17833_),
    .Y(_17834_));
 sky130_fd_sc_hd__a211o_2 _40420_ (.A1(_17741_),
    .A2(_17737_),
    .B1(_17833_),
    .C1(_17735_),
    .X(_17835_));
 sky130_fd_sc_hd__nand2_1 _40421_ (.A(_17834_),
    .B(_17835_),
    .Y(_17836_));
 sky130_fd_sc_hd__and2_1 _40422_ (.A(_17836_),
    .B(_17594_),
    .X(_17837_));
 sky130_fd_sc_hd__nor2_2 _40423_ (.A(_17765_),
    .B(_17836_),
    .Y(_17838_));
 sky130_fd_sc_hd__nor2_1 _40424_ (.A(_17717_),
    .B(_17716_),
    .Y(_17839_));
 sky130_fd_sc_hd__o21ai_2 _40425_ (.A1(_17721_),
    .A2(_17839_),
    .B1(_17718_),
    .Y(_17840_));
 sky130_fd_sc_hd__a21o_1 _40426_ (.A1(_17574_),
    .A2(_17575_),
    .B1(_17840_),
    .X(_17841_));
 sky130_fd_sc_hd__nand2_2 _40427_ (.A(_17840_),
    .B(_17576_),
    .Y(_17842_));
 sky130_fd_sc_hd__nor2_4 _40428_ (.A(_17736_),
    .B(_16884_),
    .Y(_17843_));
 sky130_fd_sc_hd__nor2_8 _40429_ (.A(_17579_),
    .B(_17843_),
    .Y(_17844_));
 sky130_vsdinv _40430_ (.A(_17844_),
    .Y(_17845_));
 sky130_fd_sc_hd__a21oi_2 _40431_ (.A1(_17841_),
    .A2(_17842_),
    .B1(_17845_),
    .Y(_17846_));
 sky130_fd_sc_hd__and3_1 _40432_ (.A(_17841_),
    .B(_17845_),
    .C(_17842_),
    .X(_17847_));
 sky130_fd_sc_hd__nor2_2 _40433_ (.A(_17682_),
    .B(_17691_),
    .Y(_17848_));
 sky130_fd_sc_hd__a21oi_4 _40434_ (.A1(_17692_),
    .A2(_17702_),
    .B1(_17848_),
    .Y(_17849_));
 sky130_fd_sc_hd__o21a_2 _40435_ (.A1(_17684_),
    .A2(_17687_),
    .B1(_17685_),
    .X(_17850_));
 sky130_vsdinv _40436_ (.A(_17850_),
    .Y(_17851_));
 sky130_fd_sc_hd__nand2_2 _40437_ (.A(_16107_),
    .B(_20084_),
    .Y(_17852_));
 sky130_fd_sc_hd__or4_4 _40438_ (.A(_13456_),
    .B(_16448_),
    .C(_16102_),
    .D(_12307_),
    .X(_17853_));
 sky130_fd_sc_hd__a22o_1 _40439_ (.A1(_15907_),
    .A2(_20088_),
    .B1(_11941_),
    .B2(_15908_),
    .X(_17854_));
 sky130_fd_sc_hd__nand2_2 _40440_ (.A(_17853_),
    .B(_17854_),
    .Y(_17855_));
 sky130_fd_sc_hd__or2_4 _40441_ (.A(_17852_),
    .B(_17855_),
    .X(_17856_));
 sky130_fd_sc_hd__nand2_4 _40442_ (.A(_17855_),
    .B(_17852_),
    .Y(_17857_));
 sky130_fd_sc_hd__nand3_4 _40443_ (.A(_17851_),
    .B(_17856_),
    .C(_17857_),
    .Y(_17858_));
 sky130_fd_sc_hd__nand2_2 _40444_ (.A(_17856_),
    .B(_17857_),
    .Y(_17859_));
 sky130_fd_sc_hd__nand2_4 _40445_ (.A(_17859_),
    .B(_17850_),
    .Y(_17860_));
 sky130_fd_sc_hd__nand2_1 _40446_ (.A(_15897_),
    .B(_10779_),
    .Y(_17861_));
 sky130_fd_sc_hd__a22o_1 _40447_ (.A1(_15924_),
    .A2(_20079_),
    .B1(_15925_),
    .B2(_20074_),
    .X(_17862_));
 sky130_fd_sc_hd__o21ai_1 _40448_ (.A1(_10988_),
    .A2(_16281_),
    .B1(_17862_),
    .Y(_17863_));
 sky130_fd_sc_hd__or2_2 _40449_ (.A(_17861_),
    .B(_17863_),
    .X(_17864_));
 sky130_fd_sc_hd__nand2_1 _40450_ (.A(_17863_),
    .B(_17861_),
    .Y(_17865_));
 sky130_fd_sc_hd__nand2_4 _40451_ (.A(_17864_),
    .B(_17865_),
    .Y(_17866_));
 sky130_fd_sc_hd__nand3_4 _40452_ (.A(_17858_),
    .B(_17860_),
    .C(_17866_),
    .Y(_17867_));
 sky130_fd_sc_hd__nand2_2 _40453_ (.A(_17859_),
    .B(_17851_),
    .Y(_17868_));
 sky130_fd_sc_hd__nand3_4 _40454_ (.A(_17856_),
    .B(_17850_),
    .C(_17857_),
    .Y(_17869_));
 sky130_vsdinv _40455_ (.A(_17866_),
    .Y(_17870_));
 sky130_fd_sc_hd__nand3_4 _40456_ (.A(_17868_),
    .B(_17869_),
    .C(_17870_),
    .Y(_17871_));
 sky130_fd_sc_hd__nand3_4 _40457_ (.A(_17849_),
    .B(_17867_),
    .C(_17871_),
    .Y(_17872_));
 sky130_fd_sc_hd__a21oi_1 _40458_ (.A1(_17688_),
    .A2(_17689_),
    .B1(_17683_),
    .Y(_17873_));
 sky130_fd_sc_hd__o21ai_2 _40459_ (.A1(_17698_),
    .A2(_17873_),
    .B1(_17690_),
    .Y(_17874_));
 sky130_fd_sc_hd__nand3_2 _40460_ (.A(_17858_),
    .B(_17860_),
    .C(_17870_),
    .Y(_17875_));
 sky130_fd_sc_hd__nand3_2 _40461_ (.A(_17868_),
    .B(_17869_),
    .C(_17866_),
    .Y(_17876_));
 sky130_fd_sc_hd__nand3_4 _40462_ (.A(_17874_),
    .B(_17875_),
    .C(_17876_),
    .Y(_17877_));
 sky130_fd_sc_hd__nand2_1 _40463_ (.A(_17714_),
    .B(_17711_),
    .Y(_17878_));
 sky130_vsdinv _40464_ (.A(_17878_),
    .Y(_17879_));
 sky130_fd_sc_hd__o21ai_4 _40465_ (.A1(_16327_),
    .A2(_16056_),
    .B1(_17696_),
    .Y(_17880_));
 sky130_fd_sc_hd__nand2_4 _40466_ (.A(net503),
    .B(_10552_),
    .Y(_17881_));
 sky130_fd_sc_hd__or2_1 _40467_ (.A(_17710_),
    .B(_17881_),
    .X(_17882_));
 sky130_fd_sc_hd__nand2_1 _40468_ (.A(_17710_),
    .B(_17881_),
    .Y(_17883_));
 sky130_fd_sc_hd__nand2_1 _40469_ (.A(_17882_),
    .B(_17883_),
    .Y(_17884_));
 sky130_fd_sc_hd__nor2_2 _40470_ (.A(_17709_),
    .B(_17884_),
    .Y(_17885_));
 sky130_fd_sc_hd__and2_1 _40471_ (.A(_17884_),
    .B(_17709_),
    .X(_17886_));
 sky130_fd_sc_hd__nor2_4 _40472_ (.A(_17885_),
    .B(_17886_),
    .Y(_17887_));
 sky130_fd_sc_hd__or2_1 _40473_ (.A(_17880_),
    .B(_17887_),
    .X(_17888_));
 sky130_fd_sc_hd__nand2_2 _40474_ (.A(_17887_),
    .B(_17880_),
    .Y(_17889_));
 sky130_fd_sc_hd__nand2_2 _40475_ (.A(_17888_),
    .B(_17889_),
    .Y(_17890_));
 sky130_fd_sc_hd__nor2_2 _40476_ (.A(_17879_),
    .B(_17890_),
    .Y(_17891_));
 sky130_fd_sc_hd__and2_1 _40477_ (.A(_17890_),
    .B(_17879_),
    .X(_17892_));
 sky130_fd_sc_hd__o2bb2ai_4 _40478_ (.A1_N(_17872_),
    .A2_N(_17877_),
    .B1(_17891_),
    .B2(_17892_),
    .Y(_17893_));
 sky130_fd_sc_hd__nand2_1 _40479_ (.A(_17890_),
    .B(_17878_),
    .Y(_17894_));
 sky130_fd_sc_hd__nand3_1 _40480_ (.A(_17879_),
    .B(_17888_),
    .C(_17889_),
    .Y(_17895_));
 sky130_fd_sc_hd__nand2_2 _40481_ (.A(_17894_),
    .B(_17895_),
    .Y(_17896_));
 sky130_fd_sc_hd__nand3_4 _40482_ (.A(_17877_),
    .B(_17872_),
    .C(_17896_),
    .Y(_17897_));
 sky130_fd_sc_hd__o21ai_1 _40483_ (.A1(_17722_),
    .A2(_17724_),
    .B1(_17704_),
    .Y(_17898_));
 sky130_fd_sc_hd__nand2_2 _40484_ (.A(_17898_),
    .B(_17708_),
    .Y(_17899_));
 sky130_fd_sc_hd__a21oi_4 _40485_ (.A1(_17893_),
    .A2(_17897_),
    .B1(_17899_),
    .Y(_17900_));
 sky130_fd_sc_hd__nand2_1 _40486_ (.A(_17706_),
    .B(_17707_),
    .Y(_17901_));
 sky130_fd_sc_hd__nor2_1 _40487_ (.A(_17681_),
    .B(_17901_),
    .Y(_17902_));
 sky130_fd_sc_hd__a2bb2oi_1 _40488_ (.A1_N(_17722_),
    .A2_N(_17724_),
    .B1(_17681_),
    .B2(_17901_),
    .Y(_17903_));
 sky130_fd_sc_hd__o211a_1 _40489_ (.A1(_17902_),
    .A2(_17903_),
    .B1(_17897_),
    .C1(_17893_),
    .X(_17904_));
 sky130_fd_sc_hd__o22ai_4 _40490_ (.A1(_17846_),
    .A2(_17847_),
    .B1(_17900_),
    .B2(_17904_),
    .Y(_17905_));
 sky130_fd_sc_hd__clkbuf_2 _40491_ (.A(_17576_),
    .X(_17906_));
 sky130_fd_sc_hd__nor2_1 _40492_ (.A(_17906_),
    .B(_17840_),
    .Y(_17907_));
 sky130_fd_sc_hd__and2_1 _40493_ (.A(_17840_),
    .B(_17906_),
    .X(_17908_));
 sky130_fd_sc_hd__o21ai_1 _40494_ (.A1(_17907_),
    .A2(_17908_),
    .B1(_17844_),
    .Y(_17909_));
 sky130_fd_sc_hd__nand3_2 _40495_ (.A(_17841_),
    .B(_17845_),
    .C(_17842_),
    .Y(_17910_));
 sky130_fd_sc_hd__nand2_2 _40496_ (.A(_17909_),
    .B(_17910_),
    .Y(_17911_));
 sky130_fd_sc_hd__nand2_1 _40497_ (.A(_17893_),
    .B(_17897_),
    .Y(_17912_));
 sky130_fd_sc_hd__nor2_1 _40498_ (.A(_17902_),
    .B(_17903_),
    .Y(_17913_));
 sky130_fd_sc_hd__nand2_1 _40499_ (.A(_17912_),
    .B(_17913_),
    .Y(_17914_));
 sky130_fd_sc_hd__nand3_4 _40500_ (.A(_17893_),
    .B(_17899_),
    .C(_17897_),
    .Y(_17915_));
 sky130_fd_sc_hd__nand3b_4 _40501_ (.A_N(_17911_),
    .B(_17914_),
    .C(_17915_),
    .Y(_17916_));
 sky130_fd_sc_hd__nand2_2 _40502_ (.A(_17749_),
    .B(_17734_),
    .Y(_17917_));
 sky130_fd_sc_hd__a21oi_4 _40503_ (.A1(_17905_),
    .A2(_17916_),
    .B1(_17917_),
    .Y(_17918_));
 sky130_vsdinv _40504_ (.A(_17734_),
    .Y(_17919_));
 sky130_fd_sc_hd__o21a_1 _40505_ (.A1(_17753_),
    .A2(_17755_),
    .B1(_17730_),
    .X(_17920_));
 sky130_fd_sc_hd__o211a_1 _40506_ (.A1(_17919_),
    .A2(_17920_),
    .B1(_17916_),
    .C1(_17905_),
    .X(_17921_));
 sky130_fd_sc_hd__o22ai_4 _40507_ (.A1(_17837_),
    .A2(_17838_),
    .B1(_17918_),
    .B2(_17921_),
    .Y(_17922_));
 sky130_fd_sc_hd__a21boi_4 _40508_ (.A1(_17758_),
    .A2(_17778_),
    .B1_N(_17750_),
    .Y(_17923_));
 sky130_fd_sc_hd__a21o_2 _40509_ (.A1(_17905_),
    .A2(_17916_),
    .B1(_17917_),
    .X(_17924_));
 sky130_fd_sc_hd__nand3_4 _40510_ (.A(_17917_),
    .B(_17905_),
    .C(_17916_),
    .Y(_17925_));
 sky130_fd_sc_hd__nand2_1 _40511_ (.A(_17836_),
    .B(_17759_),
    .Y(_17926_));
 sky130_fd_sc_hd__nand3_4 _40512_ (.A(_17834_),
    .B(_17835_),
    .C(_17594_),
    .Y(_17927_));
 sky130_fd_sc_hd__nand2_4 _40513_ (.A(_17926_),
    .B(_17927_),
    .Y(_17928_));
 sky130_fd_sc_hd__nand3_4 _40514_ (.A(_17924_),
    .B(_17925_),
    .C(_17928_),
    .Y(_17929_));
 sky130_fd_sc_hd__nand3_4 _40515_ (.A(_17922_),
    .B(_17923_),
    .C(_17929_),
    .Y(_17930_));
 sky130_fd_sc_hd__o21ai_2 _40516_ (.A1(_17918_),
    .A2(_17921_),
    .B1(_17928_),
    .Y(_17931_));
 sky130_fd_sc_hd__a21oi_2 _40517_ (.A1(_17743_),
    .A2(_17749_),
    .B1(_17748_),
    .Y(_17932_));
 sky130_fd_sc_hd__o21ai_2 _40518_ (.A1(_17770_),
    .A2(_17932_),
    .B1(_17750_),
    .Y(_17933_));
 sky130_vsdinv _40519_ (.A(_17928_),
    .Y(_17934_));
 sky130_fd_sc_hd__nand3_4 _40520_ (.A(_17924_),
    .B(_17925_),
    .C(_17934_),
    .Y(_17935_));
 sky130_fd_sc_hd__nand3_4 _40521_ (.A(_17931_),
    .B(_17933_),
    .C(_17935_),
    .Y(_17936_));
 sky130_fd_sc_hd__nand2_1 _40522_ (.A(_17769_),
    .B(_17760_),
    .Y(_17937_));
 sky130_fd_sc_hd__nand2_1 _40523_ (.A(_17937_),
    .B(_17613_),
    .Y(_17938_));
 sky130_fd_sc_hd__a21boi_2 _40524_ (.A1(_17594_),
    .A2(_17761_),
    .B1_N(_17760_),
    .Y(_17939_));
 sky130_fd_sc_hd__nand2_1 _40525_ (.A(_17939_),
    .B(_16971_),
    .Y(_17940_));
 sky130_fd_sc_hd__nand2_1 _40526_ (.A(_17938_),
    .B(_17940_),
    .Y(_17941_));
 sky130_fd_sc_hd__nor2_1 _40527_ (.A(_17796_),
    .B(_17941_),
    .Y(_17942_));
 sky130_fd_sc_hd__nor2_2 _40528_ (.A(_16971_),
    .B(_17939_),
    .Y(_17943_));
 sky130_fd_sc_hd__clkbuf_2 _40529_ (.A(_16783_),
    .X(_17944_));
 sky130_fd_sc_hd__nor2_1 _40530_ (.A(_17944_),
    .B(_17937_),
    .Y(_17945_));
 sky130_fd_sc_hd__nor2_1 _40531_ (.A(_17943_),
    .B(_17945_),
    .Y(_17946_));
 sky130_fd_sc_hd__nor2_1 _40532_ (.A(_17176_),
    .B(_17946_),
    .Y(_17947_));
 sky130_fd_sc_hd__o2bb2ai_1 _40533_ (.A1_N(_17930_),
    .A2_N(_17936_),
    .B1(_17942_),
    .B2(_17947_),
    .Y(_17948_));
 sky130_fd_sc_hd__nand2_1 _40534_ (.A(_17589_),
    .B(_17607_),
    .Y(_17949_));
 sky130_fd_sc_hd__a22oi_4 _40535_ (.A1(_17949_),
    .A2(_17593_),
    .B1(_17767_),
    .B2(_17771_),
    .Y(_17950_));
 sky130_fd_sc_hd__a21oi_4 _40536_ (.A1(_17772_),
    .A2(_17788_),
    .B1(_17950_),
    .Y(_17951_));
 sky130_fd_sc_hd__nand2_2 _40537_ (.A(_17940_),
    .B(_16592_),
    .Y(_17952_));
 sky130_fd_sc_hd__nand2_1 _40538_ (.A(_17941_),
    .B(_16982_),
    .Y(_17953_));
 sky130_fd_sc_hd__o21ai_2 _40539_ (.A1(_17943_),
    .A2(_17952_),
    .B1(_17953_),
    .Y(_17954_));
 sky130_fd_sc_hd__nand3_2 _40540_ (.A(_17936_),
    .B(_17930_),
    .C(_17954_),
    .Y(_17955_));
 sky130_fd_sc_hd__nand3_4 _40541_ (.A(_17948_),
    .B(_17951_),
    .C(_17955_),
    .Y(_17956_));
 sky130_fd_sc_hd__a31oi_4 _40542_ (.A1(_17680_),
    .A2(_17767_),
    .A3(_17771_),
    .B1(_17793_),
    .Y(_17957_));
 sky130_vsdinv _40543_ (.A(_17954_),
    .Y(_17958_));
 sky130_fd_sc_hd__nand3_2 _40544_ (.A(_17958_),
    .B(_17936_),
    .C(_17930_),
    .Y(_17959_));
 sky130_fd_sc_hd__nor2_1 _40545_ (.A(_17943_),
    .B(_17952_),
    .Y(_17960_));
 sky130_fd_sc_hd__nor2_1 _40546_ (.A(_17796_),
    .B(_17946_),
    .Y(_17961_));
 sky130_fd_sc_hd__o2bb2ai_2 _40547_ (.A1_N(_17930_),
    .A2_N(_17936_),
    .B1(_17960_),
    .B2(_17961_),
    .Y(_17962_));
 sky130_fd_sc_hd__o211ai_4 _40548_ (.A1(_17950_),
    .A2(_17957_),
    .B1(_17959_),
    .C1(_17962_),
    .Y(_17963_));
 sky130_fd_sc_hd__nand2_2 _40549_ (.A(_17785_),
    .B(_17782_),
    .Y(_17964_));
 sky130_vsdinv _40550_ (.A(_17964_),
    .Y(_17965_));
 sky130_fd_sc_hd__nor2_8 _40551_ (.A(net413),
    .B(_17965_),
    .Y(_17966_));
 sky130_fd_sc_hd__nor2_4 _40552_ (.A(_16426_),
    .B(_17964_),
    .Y(_17967_));
 sky130_fd_sc_hd__o2bb2ai_2 _40553_ (.A1_N(_17956_),
    .A2_N(_17963_),
    .B1(_17966_),
    .B2(_17967_),
    .Y(_17968_));
 sky130_fd_sc_hd__nor2_4 _40554_ (.A(_17967_),
    .B(_17966_),
    .Y(_17969_));
 sky130_fd_sc_hd__nand3_2 _40555_ (.A(_17963_),
    .B(_17956_),
    .C(_17969_),
    .Y(_17970_));
 sky130_fd_sc_hd__o211ai_4 _40556_ (.A1(_17831_),
    .A2(_17812_),
    .B1(_17968_),
    .C1(_17970_),
    .Y(_17971_));
 sky130_fd_sc_hd__a21oi_2 _40557_ (.A1(_17799_),
    .A2(_17802_),
    .B1(_17831_),
    .Y(_17972_));
 sky130_fd_sc_hd__nor2_1 _40558_ (.A(_17004_),
    .B(_17965_),
    .Y(_17973_));
 sky130_fd_sc_hd__nor2_1 _40559_ (.A(net411),
    .B(_17964_),
    .Y(_17974_));
 sky130_fd_sc_hd__o2bb2ai_1 _40560_ (.A1_N(_17956_),
    .A2_N(_17963_),
    .B1(_17973_),
    .B2(_17974_),
    .Y(_17975_));
 sky130_fd_sc_hd__nand3b_2 _40561_ (.A_N(_17969_),
    .B(_17963_),
    .C(_17956_),
    .Y(_17976_));
 sky130_fd_sc_hd__nand3_4 _40562_ (.A(_17972_),
    .B(_17975_),
    .C(_17976_),
    .Y(_17977_));
 sky130_fd_sc_hd__a21oi_1 _40563_ (.A1(_17971_),
    .A2(_17977_),
    .B1(_17810_),
    .Y(_17978_));
 sky130_fd_sc_hd__and3_1 _40564_ (.A(_17971_),
    .B(_17977_),
    .C(_17810_),
    .X(_17979_));
 sky130_fd_sc_hd__a21oi_2 _40565_ (.A1(_17804_),
    .A2(_17806_),
    .B1(_17805_),
    .Y(_17980_));
 sky130_fd_sc_hd__a21oi_1 _40566_ (.A1(_17807_),
    .A2(_17640_),
    .B1(_17980_),
    .Y(_17981_));
 sky130_fd_sc_hd__o21ai_1 _40567_ (.A1(_17978_),
    .A2(_17979_),
    .B1(_17981_),
    .Y(_17982_));
 sky130_fd_sc_hd__a31oi_2 _40568_ (.A1(_17804_),
    .A2(_17805_),
    .A3(_17806_),
    .B1(_17677_),
    .Y(_17983_));
 sky130_fd_sc_hd__a21o_1 _40569_ (.A1(_17971_),
    .A2(_17977_),
    .B1(_17810_),
    .X(_17984_));
 sky130_fd_sc_hd__nand3_1 _40570_ (.A(_17971_),
    .B(_17977_),
    .C(_17810_),
    .Y(_17985_));
 sky130_fd_sc_hd__o211ai_2 _40571_ (.A1(_17980_),
    .A2(_17983_),
    .B1(_17984_),
    .C1(_17985_),
    .Y(_17986_));
 sky130_fd_sc_hd__and2_1 _40572_ (.A(_17982_),
    .B(_17986_),
    .X(_17987_));
 sky130_fd_sc_hd__a21boi_4 _40573_ (.A1(_17827_),
    .A2(_17830_),
    .B1_N(_17987_),
    .Y(_17988_));
 sky130_fd_sc_hd__and3b_1 _40574_ (.A_N(_17987_),
    .B(_17827_),
    .C(_17830_),
    .X(_17989_));
 sky130_fd_sc_hd__nor2_4 _40575_ (.A(_17988_),
    .B(_17989_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_2 _40576_ (.A(_17910_),
    .B(_17842_),
    .Y(_17990_));
 sky130_fd_sc_hd__or2b_2 _40577_ (.A(_17990_),
    .B_N(_17320_),
    .X(_17991_));
 sky130_fd_sc_hd__nand2_2 _40578_ (.A(_17990_),
    .B(_17833_),
    .Y(_17992_));
 sky130_fd_sc_hd__a21oi_4 _40579_ (.A1(_17991_),
    .A2(_17992_),
    .B1(_17759_),
    .Y(_17993_));
 sky130_fd_sc_hd__and3_2 _40580_ (.A(_17991_),
    .B(_17759_),
    .C(_17992_),
    .X(_17994_));
 sky130_fd_sc_hd__o21ai_4 _40581_ (.A1(_17879_),
    .A2(_17890_),
    .B1(_17889_),
    .Y(_17995_));
 sky130_fd_sc_hd__and2_1 _40582_ (.A(_17995_),
    .B(_17739_),
    .X(_17996_));
 sky130_fd_sc_hd__nor2_4 _40583_ (.A(_17739_),
    .B(_17995_),
    .Y(_17997_));
 sky130_fd_sc_hd__nor2_2 _40584_ (.A(_17850_),
    .B(_17859_),
    .Y(_17998_));
 sky130_fd_sc_hd__a21oi_2 _40585_ (.A1(_17860_),
    .A2(_17870_),
    .B1(_17998_),
    .Y(_17999_));
 sky130_fd_sc_hd__nor2_1 _40586_ (.A(_10405_),
    .B(_11181_),
    .Y(_18000_));
 sky130_vsdinv _40587_ (.A(_18000_),
    .Y(_18001_));
 sky130_fd_sc_hd__or4_4 _40588_ (.A(_20088_),
    .B(_15914_),
    .C(_15916_),
    .D(_10763_),
    .X(_18002_));
 sky130_fd_sc_hd__a22o_1 _40589_ (.A1(_19831_),
    .A2(_20083_),
    .B1(_12297_),
    .B2(_18696_),
    .X(_18003_));
 sky130_fd_sc_hd__nand2_1 _40590_ (.A(_18002_),
    .B(_18003_),
    .Y(_18004_));
 sky130_fd_sc_hd__or2_4 _40591_ (.A(_18001_),
    .B(_18004_),
    .X(_18005_));
 sky130_fd_sc_hd__nand2_2 _40592_ (.A(_18004_),
    .B(_18001_),
    .Y(_18006_));
 sky130_fd_sc_hd__o21a_1 _40593_ (.A1(_17852_),
    .A2(_17855_),
    .B1(_17853_),
    .X(_18007_));
 sky130_fd_sc_hd__a21bo_1 _40594_ (.A1(_18005_),
    .A2(_18006_),
    .B1_N(_18007_),
    .X(_18008_));
 sky130_vsdinv _40595_ (.A(_18007_),
    .Y(_18009_));
 sky130_fd_sc_hd__nand3_4 _40596_ (.A(_18009_),
    .B(_18005_),
    .C(_18006_),
    .Y(_18010_));
 sky130_fd_sc_hd__nand2_4 _40597_ (.A(_18687_),
    .B(_15897_),
    .Y(_18011_));
 sky130_fd_sc_hd__and4_1 _40598_ (.A(_15924_),
    .B(_19842_),
    .C(_20070_),
    .D(_11607_),
    .X(_18012_));
 sky130_fd_sc_hd__o22a_1 _40599_ (.A1(_16094_),
    .A2(_16059_),
    .B1(_16095_),
    .B2(_16147_),
    .X(_18013_));
 sky130_fd_sc_hd__or3_1 _40600_ (.A(_18011_),
    .B(_18012_),
    .C(_18013_),
    .X(_18014_));
 sky130_fd_sc_hd__o21ai_1 _40601_ (.A1(_18012_),
    .A2(_18013_),
    .B1(_18011_),
    .Y(_18015_));
 sky130_fd_sc_hd__nand2_2 _40602_ (.A(_18014_),
    .B(_18015_),
    .Y(_18016_));
 sky130_fd_sc_hd__nand3_2 _40603_ (.A(_18008_),
    .B(_18010_),
    .C(_18016_),
    .Y(_18017_));
 sky130_fd_sc_hd__a21o_1 _40604_ (.A1(_18005_),
    .A2(_18006_),
    .B1(_18007_),
    .X(_18018_));
 sky130_fd_sc_hd__nand3_2 _40605_ (.A(_18005_),
    .B(_18007_),
    .C(_18006_),
    .Y(_18019_));
 sky130_vsdinv _40606_ (.A(_18016_),
    .Y(_18020_));
 sky130_fd_sc_hd__nand3_2 _40607_ (.A(_18018_),
    .B(_18019_),
    .C(_18020_),
    .Y(_18021_));
 sky130_fd_sc_hd__nand3_4 _40608_ (.A(_17999_),
    .B(_18017_),
    .C(_18021_),
    .Y(_18022_));
 sky130_fd_sc_hd__a21o_1 _40609_ (.A1(_17860_),
    .A2(_17870_),
    .B1(_17998_),
    .X(_18023_));
 sky130_fd_sc_hd__nand3_4 _40610_ (.A(_18008_),
    .B(_18010_),
    .C(_18020_),
    .Y(_18024_));
 sky130_fd_sc_hd__nand3_2 _40611_ (.A(_18018_),
    .B(_18019_),
    .C(_18016_),
    .Y(_18025_));
 sky130_fd_sc_hd__nand3_4 _40612_ (.A(_18023_),
    .B(_18024_),
    .C(_18025_),
    .Y(_18026_));
 sky130_vsdinv _40613_ (.A(_17882_),
    .Y(_18027_));
 sky130_fd_sc_hd__nor2_1 _40614_ (.A(_18027_),
    .B(_17885_),
    .Y(_18028_));
 sky130_fd_sc_hd__clkbuf_2 _40615_ (.A(_18028_),
    .X(_18029_));
 sky130_fd_sc_hd__buf_2 _40616_ (.A(_18029_),
    .X(_18030_));
 sky130_fd_sc_hd__o21ai_4 _40617_ (.A1(_16327_),
    .A2(_16281_),
    .B1(_17864_),
    .Y(_18031_));
 sky130_fd_sc_hd__or2_1 _40618_ (.A(_18031_),
    .B(_17887_),
    .X(_18032_));
 sky130_fd_sc_hd__clkbuf_2 _40619_ (.A(_17887_),
    .X(_18033_));
 sky130_fd_sc_hd__nand2_2 _40620_ (.A(_18033_),
    .B(_18031_),
    .Y(_18034_));
 sky130_fd_sc_hd__nand2_4 _40621_ (.A(_18032_),
    .B(_18034_),
    .Y(_18035_));
 sky130_fd_sc_hd__nor2_4 _40622_ (.A(_18030_),
    .B(_18035_),
    .Y(_18036_));
 sky130_vsdinv _40623_ (.A(_18029_),
    .Y(_18037_));
 sky130_vsdinv _40624_ (.A(_18035_),
    .Y(_18038_));
 sky130_fd_sc_hd__nor2_4 _40625_ (.A(_18037_),
    .B(_18038_),
    .Y(_18039_));
 sky130_fd_sc_hd__o2bb2ai_2 _40626_ (.A1_N(_18022_),
    .A2_N(_18026_),
    .B1(_18036_),
    .B2(_18039_),
    .Y(_18040_));
 sky130_fd_sc_hd__nor2_2 _40627_ (.A(_18037_),
    .B(_18035_),
    .Y(_18041_));
 sky130_fd_sc_hd__nor2_2 _40628_ (.A(_18030_),
    .B(_18038_),
    .Y(_18042_));
 sky130_fd_sc_hd__o211ai_4 _40629_ (.A1(_18041_),
    .A2(_18042_),
    .B1(_18022_),
    .C1(_18026_),
    .Y(_18043_));
 sky130_fd_sc_hd__nand2_2 _40630_ (.A(_17897_),
    .B(_17877_),
    .Y(_18044_));
 sky130_fd_sc_hd__a21oi_2 _40631_ (.A1(_18040_),
    .A2(_18043_),
    .B1(_18044_),
    .Y(_18045_));
 sky130_fd_sc_hd__a21oi_4 _40632_ (.A1(_17867_),
    .A2(_17871_),
    .B1(_17849_),
    .Y(_18046_));
 sky130_fd_sc_hd__a21oi_4 _40633_ (.A1(_17872_),
    .A2(_17896_),
    .B1(_18046_),
    .Y(_18047_));
 sky130_fd_sc_hd__a2bb2oi_4 _40634_ (.A1_N(_18036_),
    .A2_N(_18039_),
    .B1(_18022_),
    .B2(_18026_),
    .Y(_18048_));
 sky130_fd_sc_hd__o211a_1 _40635_ (.A1(_18041_),
    .A2(_18042_),
    .B1(_18022_),
    .C1(_18026_),
    .X(_18049_));
 sky130_fd_sc_hd__nor3_4 _40636_ (.A(_18047_),
    .B(_18048_),
    .C(_18049_),
    .Y(_18050_));
 sky130_fd_sc_hd__o22ai_4 _40637_ (.A1(_17996_),
    .A2(_17997_),
    .B1(_18045_),
    .B2(_18050_),
    .Y(_18051_));
 sky130_fd_sc_hd__o21ai_2 _40638_ (.A1(_18048_),
    .A2(_18049_),
    .B1(_18047_),
    .Y(_18052_));
 sky130_fd_sc_hd__nor2_2 _40639_ (.A(_17997_),
    .B(_17996_),
    .Y(_18053_));
 sky130_fd_sc_hd__nand3_4 _40640_ (.A(_18044_),
    .B(_18040_),
    .C(_18043_),
    .Y(_18054_));
 sky130_fd_sc_hd__nand3_4 _40641_ (.A(_18052_),
    .B(_18053_),
    .C(_18054_),
    .Y(_18055_));
 sky130_fd_sc_hd__o21ai_4 _40642_ (.A1(_17911_),
    .A2(_17900_),
    .B1(_17915_),
    .Y(_18056_));
 sky130_fd_sc_hd__a21oi_4 _40643_ (.A1(_18051_),
    .A2(_18055_),
    .B1(_18056_),
    .Y(_18057_));
 sky130_fd_sc_hd__a21oi_1 _40644_ (.A1(_17912_),
    .A2(_17913_),
    .B1(_17911_),
    .Y(_18058_));
 sky130_fd_sc_hd__o211a_2 _40645_ (.A1(_17904_),
    .A2(_18058_),
    .B1(_18055_),
    .C1(_18051_),
    .X(_18059_));
 sky130_fd_sc_hd__o22ai_4 _40646_ (.A1(_17993_),
    .A2(_17994_),
    .B1(_18057_),
    .B2(_18059_),
    .Y(_18060_));
 sky130_fd_sc_hd__nand2_1 _40647_ (.A(_17925_),
    .B(_17928_),
    .Y(_18061_));
 sky130_fd_sc_hd__nand2_1 _40648_ (.A(_18061_),
    .B(_17924_),
    .Y(_18062_));
 sky130_fd_sc_hd__a21o_1 _40649_ (.A1(_18051_),
    .A2(_18055_),
    .B1(_18056_),
    .X(_18063_));
 sky130_fd_sc_hd__and2_1 _40650_ (.A(_17990_),
    .B(_17833_),
    .X(_18064_));
 sky130_fd_sc_hd__nand2_1 _40651_ (.A(_17991_),
    .B(_17594_),
    .Y(_18065_));
 sky130_fd_sc_hd__nor2_1 _40652_ (.A(_17833_),
    .B(_17990_),
    .Y(_18066_));
 sky130_fd_sc_hd__o21ai_1 _40653_ (.A1(_18066_),
    .A2(_18064_),
    .B1(_17759_),
    .Y(_18067_));
 sky130_fd_sc_hd__o21ai_2 _40654_ (.A1(_18064_),
    .A2(_18065_),
    .B1(_18067_),
    .Y(_18068_));
 sky130_fd_sc_hd__nand3_4 _40655_ (.A(_18051_),
    .B(_18056_),
    .C(_18055_),
    .Y(_18069_));
 sky130_fd_sc_hd__nand3_2 _40656_ (.A(_18063_),
    .B(_18068_),
    .C(_18069_),
    .Y(_18070_));
 sky130_fd_sc_hd__nand3_4 _40657_ (.A(_18060_),
    .B(_18062_),
    .C(_18070_),
    .Y(_18071_));
 sky130_fd_sc_hd__o21ai_2 _40658_ (.A1(_18057_),
    .A2(_18059_),
    .B1(_18068_),
    .Y(_18072_));
 sky130_fd_sc_hd__o21ai_2 _40659_ (.A1(_17928_),
    .A2(_17918_),
    .B1(_17925_),
    .Y(_18073_));
 sky130_fd_sc_hd__o211ai_4 _40660_ (.A1(_17993_),
    .A2(_17994_),
    .B1(_18069_),
    .C1(_18063_),
    .Y(_18074_));
 sky130_fd_sc_hd__nand3_4 _40661_ (.A(_18072_),
    .B(_18073_),
    .C(_18074_),
    .Y(_18075_));
 sky130_fd_sc_hd__nand2_1 _40662_ (.A(_17927_),
    .B(_17834_),
    .Y(_18076_));
 sky130_vsdinv _40663_ (.A(_18076_),
    .Y(_18077_));
 sky130_fd_sc_hd__nand2_2 _40664_ (.A(_18077_),
    .B(_16971_),
    .Y(_18078_));
 sky130_fd_sc_hd__nand2_2 _40665_ (.A(_18076_),
    .B(_17613_),
    .Y(_18079_));
 sky130_fd_sc_hd__and3_1 _40666_ (.A(_18078_),
    .B(_16975_),
    .C(_18079_),
    .X(_18080_));
 sky130_fd_sc_hd__a21oi_4 _40667_ (.A1(_18078_),
    .A2(_18079_),
    .B1(_16975_),
    .Y(_18081_));
 sky130_fd_sc_hd__o2bb2ai_4 _40668_ (.A1_N(_18071_),
    .A2_N(_18075_),
    .B1(_18080_),
    .B2(_18081_),
    .Y(_18082_));
 sky130_fd_sc_hd__nor2_2 _40669_ (.A(_18081_),
    .B(_18080_),
    .Y(_18083_));
 sky130_fd_sc_hd__nand3_4 _40670_ (.A(_18083_),
    .B(_18075_),
    .C(_18071_),
    .Y(_18084_));
 sky130_vsdinv _40671_ (.A(_17935_),
    .Y(_18085_));
 sky130_fd_sc_hd__nand2_1 _40672_ (.A(_17931_),
    .B(_17933_),
    .Y(_18086_));
 sky130_fd_sc_hd__o2bb2ai_4 _40673_ (.A1_N(_17930_),
    .A2_N(_17958_),
    .B1(_18085_),
    .B2(_18086_),
    .Y(_18087_));
 sky130_fd_sc_hd__a21oi_4 _40674_ (.A1(_18082_),
    .A2(_18084_),
    .B1(_18087_),
    .Y(_18088_));
 sky130_fd_sc_hd__a31oi_1 _40675_ (.A1(_17922_),
    .A2(_17923_),
    .A3(_17929_),
    .B1(_17954_),
    .Y(_18089_));
 sky130_vsdinv _40676_ (.A(_17936_),
    .Y(_18090_));
 sky130_fd_sc_hd__o211a_1 _40677_ (.A1(_18089_),
    .A2(_18090_),
    .B1(_18084_),
    .C1(_18082_),
    .X(_18091_));
 sky130_fd_sc_hd__and3_1 _40678_ (.A(_17952_),
    .B(_15754_),
    .C(_17938_),
    .X(_18092_));
 sky130_fd_sc_hd__and2_2 _40679_ (.A(_17952_),
    .B(_17938_),
    .X(_18093_));
 sky130_fd_sc_hd__nor2_8 _40680_ (.A(_14354_),
    .B(_18093_),
    .Y(_18094_));
 sky130_fd_sc_hd__or2_2 _40681_ (.A(_18092_),
    .B(_18094_),
    .X(_18095_));
 sky130_vsdinv _40682_ (.A(_18095_),
    .Y(_18096_));
 sky130_fd_sc_hd__o21ai_2 _40683_ (.A1(_18088_),
    .A2(_18091_),
    .B1(_18096_),
    .Y(_18097_));
 sky130_fd_sc_hd__a21boi_2 _40684_ (.A1(_17956_),
    .A2(_17969_),
    .B1_N(_17963_),
    .Y(_18098_));
 sky130_fd_sc_hd__a21o_1 _40685_ (.A1(_18082_),
    .A2(_18084_),
    .B1(_18087_),
    .X(_18099_));
 sky130_fd_sc_hd__nand3_4 _40686_ (.A(_18087_),
    .B(_18082_),
    .C(_18084_),
    .Y(_18100_));
 sky130_fd_sc_hd__nand3_2 _40687_ (.A(_18099_),
    .B(_18100_),
    .C(_18095_),
    .Y(_18101_));
 sky130_fd_sc_hd__nand3_4 _40688_ (.A(_18097_),
    .B(_18098_),
    .C(_18101_),
    .Y(_18102_));
 sky130_fd_sc_hd__o22ai_4 _40689_ (.A1(_18094_),
    .A2(_18092_),
    .B1(_18088_),
    .B2(_18091_),
    .Y(_18103_));
 sky130_fd_sc_hd__nand2_1 _40690_ (.A(_17956_),
    .B(_17969_),
    .Y(_18104_));
 sky130_fd_sc_hd__nand2_1 _40691_ (.A(_18104_),
    .B(_17963_),
    .Y(_18105_));
 sky130_fd_sc_hd__nand3_2 _40692_ (.A(_18099_),
    .B(_18100_),
    .C(_18096_),
    .Y(_18106_));
 sky130_fd_sc_hd__nand3_4 _40693_ (.A(_18103_),
    .B(_18105_),
    .C(_18106_),
    .Y(_18107_));
 sky130_fd_sc_hd__a21oi_1 _40694_ (.A1(_18102_),
    .A2(_18107_),
    .B1(_17966_),
    .Y(_18108_));
 sky130_fd_sc_hd__and3_1 _40695_ (.A(_18102_),
    .B(_18107_),
    .C(_17966_),
    .X(_18109_));
 sky130_fd_sc_hd__nand2_1 _40696_ (.A(_17977_),
    .B(_17810_),
    .Y(_18110_));
 sky130_fd_sc_hd__nand2_1 _40697_ (.A(_18110_),
    .B(_17971_),
    .Y(_18111_));
 sky130_fd_sc_hd__o21bai_1 _40698_ (.A1(_18108_),
    .A2(_18109_),
    .B1_N(_18111_),
    .Y(_18112_));
 sky130_fd_sc_hd__a21o_1 _40699_ (.A1(_18102_),
    .A2(_18107_),
    .B1(_17966_),
    .X(_18113_));
 sky130_fd_sc_hd__nand3_2 _40700_ (.A(_18102_),
    .B(_18107_),
    .C(_17966_),
    .Y(_18114_));
 sky130_fd_sc_hd__nand3_2 _40701_ (.A(_18113_),
    .B(_18114_),
    .C(_18111_),
    .Y(_18115_));
 sky130_fd_sc_hd__and2_1 _40702_ (.A(_18112_),
    .B(_18115_),
    .X(_18116_));
 sky130_fd_sc_hd__nand2_1 _40703_ (.A(_18116_),
    .B(_17986_),
    .Y(_18117_));
 sky130_vsdinv _40704_ (.A(_17986_),
    .Y(_18118_));
 sky130_fd_sc_hd__o21bai_2 _40705_ (.A1(_18118_),
    .A2(_17988_),
    .B1_N(_18116_),
    .Y(_18119_));
 sky130_fd_sc_hd__o21ai_4 _40706_ (.A1(_17988_),
    .A2(_18117_),
    .B1(_18119_),
    .Y(_02678_));
 sky130_fd_sc_hd__o21ai_4 _40707_ (.A1(_18095_),
    .A2(_18088_),
    .B1(_18100_),
    .Y(_18120_));
 sky130_fd_sc_hd__nor2_1 _40708_ (.A(_13024_),
    .B(_16095_),
    .Y(_18121_));
 sky130_fd_sc_hd__a21oi_2 _40709_ (.A1(_19837_),
    .A2(_20071_),
    .B1(_18121_),
    .Y(_18122_));
 sky130_fd_sc_hd__and3_1 _40710_ (.A(_18121_),
    .B(_19837_),
    .C(_10779_),
    .X(_18123_));
 sky130_fd_sc_hd__nor2_4 _40711_ (.A(_18122_),
    .B(_18123_),
    .Y(_18124_));
 sky130_fd_sc_hd__xnor2_4 _40712_ (.A(_18011_),
    .B(_18124_),
    .Y(_18125_));
 sky130_fd_sc_hd__nand2_1 _40713_ (.A(_19834_),
    .B(_20075_),
    .Y(_18126_));
 sky130_fd_sc_hd__or4_4 _40714_ (.A(_20083_),
    .B(_16448_),
    .C(_15916_),
    .D(_11181_),
    .X(_18127_));
 sky130_fd_sc_hd__a22o_1 _40715_ (.A1(_19831_),
    .A2(_13647_),
    .B1(_10763_),
    .B2(_15908_),
    .X(_18128_));
 sky130_fd_sc_hd__nand2_1 _40716_ (.A(_18127_),
    .B(_18128_),
    .Y(_18129_));
 sky130_fd_sc_hd__or2_2 _40717_ (.A(_18126_),
    .B(_18129_),
    .X(_18130_));
 sky130_fd_sc_hd__nand2_1 _40718_ (.A(_18129_),
    .B(_18126_),
    .Y(_18131_));
 sky130_fd_sc_hd__nand2_2 _40719_ (.A(_18130_),
    .B(_18131_),
    .Y(_18132_));
 sky130_fd_sc_hd__a21o_1 _40720_ (.A1(_18002_),
    .A2(_18005_),
    .B1(_18132_),
    .X(_18133_));
 sky130_fd_sc_hd__nand3_4 _40721_ (.A(_18132_),
    .B(_18002_),
    .C(_18005_),
    .Y(_18134_));
 sky130_fd_sc_hd__nand2_1 _40722_ (.A(_18133_),
    .B(_18134_),
    .Y(_18135_));
 sky130_fd_sc_hd__nor2_2 _40723_ (.A(_18125_),
    .B(_18135_),
    .Y(_18136_));
 sky130_fd_sc_hd__and2_1 _40724_ (.A(_18135_),
    .B(_18125_),
    .X(_18137_));
 sky130_fd_sc_hd__and2_1 _40725_ (.A(_18024_),
    .B(_18010_),
    .X(_18138_));
 sky130_fd_sc_hd__o21bai_4 _40726_ (.A1(_18136_),
    .A2(_18137_),
    .B1_N(_18138_),
    .Y(_18139_));
 sky130_fd_sc_hd__nand2_1 _40727_ (.A(_18135_),
    .B(_18125_),
    .Y(_18140_));
 sky130_fd_sc_hd__nand3b_4 _40728_ (.A_N(_18136_),
    .B(_18138_),
    .C(_18140_),
    .Y(_18141_));
 sky130_fd_sc_hd__o21bai_2 _40729_ (.A1(_18011_),
    .A2(_18013_),
    .B1_N(_18012_),
    .Y(_18142_));
 sky130_fd_sc_hd__or2_1 _40730_ (.A(_18142_),
    .B(_17887_),
    .X(_18143_));
 sky130_fd_sc_hd__nand2_1 _40731_ (.A(_18033_),
    .B(_18142_),
    .Y(_18144_));
 sky130_fd_sc_hd__nand2_1 _40732_ (.A(_18143_),
    .B(_18144_),
    .Y(_18145_));
 sky130_fd_sc_hd__or2_1 _40733_ (.A(_18028_),
    .B(_18145_),
    .X(_18146_));
 sky130_fd_sc_hd__nand2_1 _40734_ (.A(_18145_),
    .B(_18029_),
    .Y(_18147_));
 sky130_fd_sc_hd__and2_2 _40735_ (.A(_18146_),
    .B(_18147_),
    .X(_18148_));
 sky130_fd_sc_hd__a21o_1 _40736_ (.A1(_18139_),
    .A2(_18141_),
    .B1(_18148_),
    .X(_18149_));
 sky130_fd_sc_hd__nand3_4 _40737_ (.A(_18139_),
    .B(_18141_),
    .C(_18148_),
    .Y(_18150_));
 sky130_fd_sc_hd__nand2_2 _40738_ (.A(_18043_),
    .B(_18026_),
    .Y(_18151_));
 sky130_fd_sc_hd__a21o_2 _40739_ (.A1(_18149_),
    .A2(_18150_),
    .B1(_18151_),
    .X(_18152_));
 sky130_fd_sc_hd__nand3_4 _40740_ (.A(_18149_),
    .B(_18150_),
    .C(_18151_),
    .Y(_18153_));
 sky130_fd_sc_hd__o21ai_2 _40741_ (.A1(_18029_),
    .A2(_18035_),
    .B1(_18034_),
    .Y(_18154_));
 sky130_fd_sc_hd__or2_1 _40742_ (.A(_17906_),
    .B(_18154_),
    .X(_18155_));
 sky130_fd_sc_hd__nand2_2 _40743_ (.A(_18154_),
    .B(_17906_),
    .Y(_18156_));
 sky130_fd_sc_hd__nand2_4 _40744_ (.A(_18155_),
    .B(_18156_),
    .Y(_18157_));
 sky130_fd_sc_hd__xor2_4 _40745_ (.A(_17844_),
    .B(_18157_),
    .X(_18158_));
 sky130_fd_sc_hd__a21o_1 _40746_ (.A1(_18152_),
    .A2(_18153_),
    .B1(_18158_),
    .X(_18159_));
 sky130_fd_sc_hd__nand2_2 _40747_ (.A(_18055_),
    .B(_18054_),
    .Y(_18160_));
 sky130_fd_sc_hd__nand3_4 _40748_ (.A(_18152_),
    .B(_18153_),
    .C(_18158_),
    .Y(_18161_));
 sky130_fd_sc_hd__nand3_4 _40749_ (.A(_18159_),
    .B(_18160_),
    .C(_18161_),
    .Y(_18162_));
 sky130_fd_sc_hd__a21oi_2 _40750_ (.A1(_18152_),
    .A2(_18153_),
    .B1(_18158_),
    .Y(_18163_));
 sky130_vsdinv _40751_ (.A(_18161_),
    .Y(_18164_));
 sky130_fd_sc_hd__o21bai_4 _40752_ (.A1(_18163_),
    .A2(_18164_),
    .B1_N(_18160_),
    .Y(_18165_));
 sky130_fd_sc_hd__a21o_1 _40753_ (.A1(_17995_),
    .A2(_17737_),
    .B1(_17735_),
    .X(_18166_));
 sky130_fd_sc_hd__nor2_1 _40754_ (.A(_17323_),
    .B(_18166_),
    .Y(_18167_));
 sky130_fd_sc_hd__and2_1 _40755_ (.A(_18166_),
    .B(_17319_),
    .X(_18168_));
 sky130_fd_sc_hd__nor2_1 _40756_ (.A(_18167_),
    .B(_18168_),
    .Y(_18169_));
 sky130_fd_sc_hd__and2_1 _40757_ (.A(_18169_),
    .B(_17393_),
    .X(_18170_));
 sky130_fd_sc_hd__nor2_2 _40758_ (.A(_17765_),
    .B(_18169_),
    .Y(_18171_));
 sky130_fd_sc_hd__o2bb2ai_4 _40759_ (.A1_N(_18162_),
    .A2_N(_18165_),
    .B1(_18170_),
    .B2(_18171_),
    .Y(_18172_));
 sky130_fd_sc_hd__or2_2 _40760_ (.A(_18171_),
    .B(_18170_),
    .X(_18173_));
 sky130_fd_sc_hd__nand3b_4 _40761_ (.A_N(_18173_),
    .B(_18165_),
    .C(_18162_),
    .Y(_18174_));
 sky130_fd_sc_hd__nor2_1 _40762_ (.A(_18057_),
    .B(_18068_),
    .Y(_18175_));
 sky130_fd_sc_hd__nor2_2 _40763_ (.A(_18059_),
    .B(_18175_),
    .Y(_18176_));
 sky130_vsdinv _40764_ (.A(_18176_),
    .Y(_18177_));
 sky130_fd_sc_hd__a21oi_4 _40765_ (.A1(_18172_),
    .A2(_18174_),
    .B1(_18177_),
    .Y(_18178_));
 sky130_fd_sc_hd__nand3_4 _40766_ (.A(_18172_),
    .B(_18174_),
    .C(_18177_),
    .Y(_18179_));
 sky130_vsdinv _40767_ (.A(_18179_),
    .Y(_18180_));
 sky130_fd_sc_hd__nand2_1 _40768_ (.A(_18065_),
    .B(_17992_),
    .Y(_18181_));
 sky130_fd_sc_hd__or2_1 _40769_ (.A(_17613_),
    .B(_18181_),
    .X(_18182_));
 sky130_fd_sc_hd__nand2_1 _40770_ (.A(_18181_),
    .B(_17944_),
    .Y(_18183_));
 sky130_fd_sc_hd__nand2_1 _40771_ (.A(_18182_),
    .B(_18183_),
    .Y(_18184_));
 sky130_fd_sc_hd__or2_2 _40772_ (.A(_17176_),
    .B(_18184_),
    .X(_18185_));
 sky130_fd_sc_hd__nand2_1 _40773_ (.A(_18184_),
    .B(_17176_),
    .Y(_18186_));
 sky130_fd_sc_hd__nand2_4 _40774_ (.A(_18185_),
    .B(_18186_),
    .Y(_18187_));
 sky130_fd_sc_hd__o21bai_2 _40775_ (.A1(_18178_),
    .A2(_18180_),
    .B1_N(_18187_),
    .Y(_18188_));
 sky130_fd_sc_hd__nand2_2 _40776_ (.A(_18084_),
    .B(_18075_),
    .Y(_18189_));
 sky130_vsdinv _40777_ (.A(_18189_),
    .Y(_18190_));
 sky130_fd_sc_hd__nand3b_4 _40778_ (.A_N(_18178_),
    .B(_18179_),
    .C(_18187_),
    .Y(_18191_));
 sky130_fd_sc_hd__nand3_4 _40779_ (.A(_18188_),
    .B(_18190_),
    .C(_18191_),
    .Y(_18192_));
 sky130_fd_sc_hd__o21ai_2 _40780_ (.A1(_18178_),
    .A2(_18180_),
    .B1(_18187_),
    .Y(_18193_));
 sky130_fd_sc_hd__nand2_1 _40781_ (.A(_18172_),
    .B(_18174_),
    .Y(_18194_));
 sky130_fd_sc_hd__a21oi_2 _40782_ (.A1(_18194_),
    .A2(_18176_),
    .B1(_18187_),
    .Y(_18195_));
 sky130_fd_sc_hd__nand2_2 _40783_ (.A(_18195_),
    .B(_18179_),
    .Y(_18196_));
 sky130_fd_sc_hd__nand3_4 _40784_ (.A(_18193_),
    .B(_18189_),
    .C(_18196_),
    .Y(_18197_));
 sky130_vsdinv _40785_ (.A(_18079_),
    .Y(_18198_));
 sky130_fd_sc_hd__and2_2 _40786_ (.A(_18078_),
    .B(_17796_),
    .X(_18199_));
 sky130_fd_sc_hd__nor2_8 _40787_ (.A(_18198_),
    .B(_18199_),
    .Y(_18200_));
 sky130_fd_sc_hd__and2_1 _40788_ (.A(_18200_),
    .B(_17004_),
    .X(_18201_));
 sky130_fd_sc_hd__nor2_2 _40789_ (.A(_17633_),
    .B(_18200_),
    .Y(_18202_));
 sky130_fd_sc_hd__o2bb2ai_2 _40790_ (.A1_N(_18192_),
    .A2_N(_18197_),
    .B1(_18201_),
    .B2(_18202_),
    .Y(_18203_));
 sky130_fd_sc_hd__nor2_2 _40791_ (.A(_18202_),
    .B(_18201_),
    .Y(_18204_));
 sky130_fd_sc_hd__nand3_2 _40792_ (.A(_18197_),
    .B(_18192_),
    .C(_18204_),
    .Y(_18205_));
 sky130_fd_sc_hd__nand3b_4 _40793_ (.A_N(_18120_),
    .B(_18203_),
    .C(_18205_),
    .Y(_18206_));
 sky130_fd_sc_hd__nor2_4 _40794_ (.A(_16818_),
    .B(_18200_),
    .Y(_18207_));
 sky130_fd_sc_hd__nand2_1 _40795_ (.A(_18200_),
    .B(_16818_),
    .Y(_18208_));
 sky130_vsdinv _40796_ (.A(_18208_),
    .Y(_18209_));
 sky130_fd_sc_hd__o2bb2ai_2 _40797_ (.A1_N(_18192_),
    .A2_N(_18197_),
    .B1(_18207_),
    .B2(_18209_),
    .Y(_18210_));
 sky130_vsdinv _40798_ (.A(_18204_),
    .Y(_18211_));
 sky130_fd_sc_hd__nand3_4 _40799_ (.A(_18197_),
    .B(_18192_),
    .C(_18211_),
    .Y(_18212_));
 sky130_fd_sc_hd__nand3_4 _40800_ (.A(_18210_),
    .B(_18120_),
    .C(_18212_),
    .Y(_18213_));
 sky130_fd_sc_hd__a21oi_4 _40801_ (.A1(_18206_),
    .A2(_18213_),
    .B1(_18094_),
    .Y(_18214_));
 sky130_fd_sc_hd__and3_1 _40802_ (.A(_18206_),
    .B(_18213_),
    .C(_18094_),
    .X(_18215_));
 sky130_fd_sc_hd__nand2_2 _40803_ (.A(_18114_),
    .B(_18107_),
    .Y(_18216_));
 sky130_fd_sc_hd__o21bai_4 _40804_ (.A1(_18214_),
    .A2(_18215_),
    .B1_N(_18216_),
    .Y(_18217_));
 sky130_fd_sc_hd__nand3_2 _40805_ (.A(_18206_),
    .B(_18213_),
    .C(_18094_),
    .Y(_18218_));
 sky130_fd_sc_hd__nand3b_4 _40806_ (.A_N(_18214_),
    .B(_18216_),
    .C(_18218_),
    .Y(_18219_));
 sky130_fd_sc_hd__nand2_1 _40807_ (.A(_18217_),
    .B(_18219_),
    .Y(_18220_));
 sky130_fd_sc_hd__and4_1 _40808_ (.A(_18112_),
    .B(_17982_),
    .C(_17986_),
    .D(_18115_),
    .X(_18221_));
 sky130_fd_sc_hd__nand2_1 _40809_ (.A(_17826_),
    .B(_18221_),
    .Y(_18222_));
 sky130_fd_sc_hd__o21bai_4 _40810_ (.A1(_17664_),
    .A2(_17673_),
    .B1_N(_18222_),
    .Y(_18223_));
 sky130_fd_sc_hd__a21bo_1 _40811_ (.A1(_18118_),
    .A2(_18112_),
    .B1_N(_18115_),
    .X(_18224_));
 sky130_fd_sc_hd__a21oi_4 _40812_ (.A1(_17829_),
    .A2(_18221_),
    .B1(_18224_),
    .Y(_18225_));
 sky130_fd_sc_hd__nand2_2 _40813_ (.A(_18223_),
    .B(_18225_),
    .Y(_18226_));
 sky130_fd_sc_hd__xnor2_2 _40814_ (.A(_18220_),
    .B(_18226_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_2 _40815_ (.A(_18185_),
    .B(_18183_),
    .Y(_18227_));
 sky130_vsdinv _40816_ (.A(_18227_),
    .Y(_18228_));
 sky130_fd_sc_hd__nor2_8 _40817_ (.A(net411),
    .B(_18228_),
    .Y(_18229_));
 sky130_fd_sc_hd__nor2_4 _40818_ (.A(_17633_),
    .B(_18227_),
    .Y(_18230_));
 sky130_fd_sc_hd__a21boi_4 _40819_ (.A1(_18148_),
    .A2(_18141_),
    .B1_N(_18139_),
    .Y(_18231_));
 sky130_fd_sc_hd__nand2_1 _40820_ (.A(_19834_),
    .B(_20071_),
    .Y(_18232_));
 sky130_fd_sc_hd__or4_4 _40821_ (.A(_20080_),
    .B(_11276_),
    .C(_16103_),
    .D(_10767_),
    .X(_18233_));
 sky130_fd_sc_hd__a22o_1 _40822_ (.A1(_19831_),
    .A2(_20075_),
    .B1(_11181_),
    .B2(_18696_),
    .X(_18234_));
 sky130_fd_sc_hd__nand2_1 _40823_ (.A(_18233_),
    .B(_18234_),
    .Y(_18235_));
 sky130_fd_sc_hd__or2_2 _40824_ (.A(_18232_),
    .B(_18235_),
    .X(_18236_));
 sky130_fd_sc_hd__nand2_1 _40825_ (.A(_18235_),
    .B(_18232_),
    .Y(_18237_));
 sky130_fd_sc_hd__nand2_2 _40826_ (.A(_18236_),
    .B(_18237_),
    .Y(_18238_));
 sky130_vsdinv _40827_ (.A(_18238_),
    .Y(_18239_));
 sky130_fd_sc_hd__nand2_1 _40828_ (.A(_18130_),
    .B(_18127_),
    .Y(_18240_));
 sky130_fd_sc_hd__nand2_2 _40829_ (.A(_18239_),
    .B(_18240_),
    .Y(_18241_));
 sky130_fd_sc_hd__and2_1 _40830_ (.A(_18130_),
    .B(_18127_),
    .X(_18242_));
 sky130_fd_sc_hd__nand2_2 _40831_ (.A(_18242_),
    .B(_18238_),
    .Y(_18243_));
 sky130_fd_sc_hd__o21ai_1 _40832_ (.A1(_19837_),
    .A2(_19842_),
    .B1(_18688_),
    .Y(_18244_));
 sky130_fd_sc_hd__and3_1 _40833_ (.A(_18688_),
    .B(_19837_),
    .C(_19842_),
    .X(_18245_));
 sky130_fd_sc_hd__nor2_1 _40834_ (.A(_18244_),
    .B(_18245_),
    .Y(_18246_));
 sky130_fd_sc_hd__nand2_2 _40835_ (.A(_18246_),
    .B(_19845_),
    .Y(_18247_));
 sky130_fd_sc_hd__o21ai_2 _40836_ (.A1(_18244_),
    .A2(_18245_),
    .B1(_18011_),
    .Y(_18248_));
 sky130_fd_sc_hd__nand2_4 _40837_ (.A(_18247_),
    .B(_18248_),
    .Y(_18249_));
 sky130_fd_sc_hd__a21o_1 _40838_ (.A1(_18241_),
    .A2(_18243_),
    .B1(_18249_),
    .X(_18250_));
 sky130_fd_sc_hd__nand3_4 _40839_ (.A(_18241_),
    .B(_18243_),
    .C(_18249_),
    .Y(_18251_));
 sky130_fd_sc_hd__a21boi_4 _40840_ (.A1(_18134_),
    .A2(_18125_),
    .B1_N(_18133_),
    .Y(_18252_));
 sky130_fd_sc_hd__a21oi_4 _40841_ (.A1(_18250_),
    .A2(_18251_),
    .B1(_18252_),
    .Y(_18253_));
 sky130_vsdinv _40842_ (.A(_18253_),
    .Y(_18254_));
 sky130_fd_sc_hd__nand3_4 _40843_ (.A(_18250_),
    .B(_18252_),
    .C(_18251_),
    .Y(_18255_));
 sky130_fd_sc_hd__a31o_1 _40844_ (.A1(_18124_),
    .A2(_18688_),
    .A3(_19845_),
    .B1(_18123_),
    .X(_18256_));
 sky130_fd_sc_hd__or2_1 _40845_ (.A(_18033_),
    .B(_18256_),
    .X(_18257_));
 sky130_fd_sc_hd__nand2_2 _40846_ (.A(_18256_),
    .B(_18033_),
    .Y(_18258_));
 sky130_fd_sc_hd__nand2_1 _40847_ (.A(_18257_),
    .B(_18258_),
    .Y(_18259_));
 sky130_fd_sc_hd__or2_2 _40848_ (.A(_18029_),
    .B(_18259_),
    .X(_18260_));
 sky130_fd_sc_hd__nand2_1 _40849_ (.A(_18259_),
    .B(_18030_),
    .Y(_18261_));
 sky130_fd_sc_hd__nand2_2 _40850_ (.A(_18260_),
    .B(_18261_),
    .Y(_18262_));
 sky130_vsdinv _40851_ (.A(_18262_),
    .Y(_18263_));
 sky130_fd_sc_hd__nand3_2 _40852_ (.A(_18254_),
    .B(_18255_),
    .C(_18263_),
    .Y(_18264_));
 sky130_vsdinv _40853_ (.A(_18255_),
    .Y(_18265_));
 sky130_fd_sc_hd__o21ai_2 _40854_ (.A1(_18253_),
    .A2(_18265_),
    .B1(_18262_),
    .Y(_18266_));
 sky130_fd_sc_hd__nand3b_4 _40855_ (.A_N(_18231_),
    .B(_18264_),
    .C(_18266_),
    .Y(_18267_));
 sky130_fd_sc_hd__nand3_2 _40856_ (.A(_18254_),
    .B(_18255_),
    .C(_18262_),
    .Y(_18268_));
 sky130_fd_sc_hd__o21ai_2 _40857_ (.A1(_18253_),
    .A2(_18265_),
    .B1(_18263_),
    .Y(_18269_));
 sky130_fd_sc_hd__nand3_4 _40858_ (.A(_18231_),
    .B(_18268_),
    .C(_18269_),
    .Y(_18270_));
 sky130_fd_sc_hd__nand2_2 _40859_ (.A(_18146_),
    .B(_18144_),
    .Y(_18271_));
 sky130_fd_sc_hd__nor2_2 _40860_ (.A(_17906_),
    .B(_18271_),
    .Y(_18272_));
 sky130_vsdinv _40861_ (.A(_18272_),
    .Y(_18273_));
 sky130_fd_sc_hd__nand2_2 _40862_ (.A(_18271_),
    .B(_17906_),
    .Y(_18274_));
 sky130_fd_sc_hd__a21oi_4 _40863_ (.A1(_18273_),
    .A2(_18274_),
    .B1(_17845_),
    .Y(_18275_));
 sky130_fd_sc_hd__and3_2 _40864_ (.A(_18273_),
    .B(_17845_),
    .C(_18274_),
    .X(_18276_));
 sky130_fd_sc_hd__nor2_8 _40865_ (.A(_18275_),
    .B(_18276_),
    .Y(_18277_));
 sky130_fd_sc_hd__a21oi_4 _40866_ (.A1(_18267_),
    .A2(_18270_),
    .B1(_18277_),
    .Y(_18278_));
 sky130_fd_sc_hd__nand2_1 _40867_ (.A(_18161_),
    .B(_18153_),
    .Y(_18279_));
 sky130_fd_sc_hd__nand3_4 _40868_ (.A(_18267_),
    .B(_18277_),
    .C(_18270_),
    .Y(_18280_));
 sky130_fd_sc_hd__nand3b_4 _40869_ (.A_N(_18278_),
    .B(_18279_),
    .C(_18280_),
    .Y(_18281_));
 sky130_fd_sc_hd__a21o_1 _40870_ (.A1(_18273_),
    .A2(_18274_),
    .B1(_17845_),
    .X(_18282_));
 sky130_fd_sc_hd__or2b_1 _40871_ (.A(_18276_),
    .B_N(_18282_),
    .X(_18283_));
 sky130_fd_sc_hd__nand2_1 _40872_ (.A(_18267_),
    .B(_18270_),
    .Y(_18284_));
 sky130_fd_sc_hd__nor2_2 _40873_ (.A(_18283_),
    .B(_18284_),
    .Y(_18285_));
 sky130_fd_sc_hd__a21boi_2 _40874_ (.A1(_18152_),
    .A2(_18158_),
    .B1_N(_18153_),
    .Y(_18286_));
 sky130_fd_sc_hd__o21ai_4 _40875_ (.A1(_18278_),
    .A2(_18285_),
    .B1(_18286_),
    .Y(_18287_));
 sky130_fd_sc_hd__o21a_1 _40876_ (.A1(_17844_),
    .A2(_18157_),
    .B1(_18156_),
    .X(_18288_));
 sky130_fd_sc_hd__nand2_2 _40877_ (.A(_18288_),
    .B(_17320_),
    .Y(_18289_));
 sky130_fd_sc_hd__o21ai_1 _40878_ (.A1(_17844_),
    .A2(_18157_),
    .B1(_18156_),
    .Y(_18290_));
 sky130_fd_sc_hd__nand2_2 _40879_ (.A(_18290_),
    .B(_17833_),
    .Y(_18291_));
 sky130_fd_sc_hd__a21oi_4 _40880_ (.A1(_18289_),
    .A2(_18291_),
    .B1(_17765_),
    .Y(_18292_));
 sky130_fd_sc_hd__and3_2 _40881_ (.A(_18289_),
    .B(_17765_),
    .C(_18291_),
    .X(_18293_));
 sky130_fd_sc_hd__o2bb2ai_4 _40882_ (.A1_N(_18281_),
    .A2_N(_18287_),
    .B1(_18292_),
    .B2(_18293_),
    .Y(_18294_));
 sky130_fd_sc_hd__nor2_8 _40883_ (.A(_18292_),
    .B(_18293_),
    .Y(_18295_));
 sky130_fd_sc_hd__nand3_4 _40884_ (.A(_18287_),
    .B(_18281_),
    .C(_18295_),
    .Y(_18296_));
 sky130_fd_sc_hd__a21oi_2 _40885_ (.A1(_18159_),
    .A2(_18161_),
    .B1(_18160_),
    .Y(_18297_));
 sky130_fd_sc_hd__o21ai_4 _40886_ (.A1(_18173_),
    .A2(_18297_),
    .B1(_18162_),
    .Y(_18298_));
 sky130_fd_sc_hd__a21oi_4 _40887_ (.A1(_18294_),
    .A2(_18296_),
    .B1(_18298_),
    .Y(_18299_));
 sky130_fd_sc_hd__and3_2 _40888_ (.A(_18294_),
    .B(_18298_),
    .C(_18296_),
    .X(_18300_));
 sky130_fd_sc_hd__or2_1 _40889_ (.A(_18168_),
    .B(_18170_),
    .X(_18301_));
 sky130_fd_sc_hd__nand2_1 _40890_ (.A(_18301_),
    .B(_17944_),
    .Y(_18302_));
 sky130_vsdinv _40891_ (.A(_18302_),
    .Y(_18303_));
 sky130_fd_sc_hd__or2_1 _40892_ (.A(_17944_),
    .B(_18301_),
    .X(_18304_));
 sky130_fd_sc_hd__nand2_2 _40893_ (.A(_18304_),
    .B(_17796_),
    .Y(_18305_));
 sky130_fd_sc_hd__nand2_1 _40894_ (.A(_18304_),
    .B(_18302_),
    .Y(_18306_));
 sky130_fd_sc_hd__nand2_2 _40895_ (.A(_18306_),
    .B(_17176_),
    .Y(_18307_));
 sky130_fd_sc_hd__o21ai_4 _40896_ (.A1(_18303_),
    .A2(_18305_),
    .B1(_18307_),
    .Y(_18308_));
 sky130_fd_sc_hd__o21ai_4 _40897_ (.A1(_18299_),
    .A2(_18300_),
    .B1(_18308_),
    .Y(_18309_));
 sky130_fd_sc_hd__a21oi_1 _40898_ (.A1(_18287_),
    .A2(_18281_),
    .B1(_18295_),
    .Y(_18310_));
 sky130_fd_sc_hd__and3_1 _40899_ (.A(_18287_),
    .B(_18281_),
    .C(_18295_),
    .X(_18311_));
 sky130_fd_sc_hd__o21bai_2 _40900_ (.A1(_18310_),
    .A2(_18311_),
    .B1_N(_18298_),
    .Y(_18312_));
 sky130_fd_sc_hd__o21a_1 _40901_ (.A1(_18303_),
    .A2(_18305_),
    .B1(_18307_),
    .X(_18313_));
 sky130_fd_sc_hd__nand3_4 _40902_ (.A(_18294_),
    .B(_18298_),
    .C(_18296_),
    .Y(_18314_));
 sky130_fd_sc_hd__nand3_4 _40903_ (.A(_18312_),
    .B(_18313_),
    .C(_18314_),
    .Y(_18315_));
 sky130_fd_sc_hd__o21ai_4 _40904_ (.A1(_18187_),
    .A2(_18178_),
    .B1(_18179_),
    .Y(_18316_));
 sky130_fd_sc_hd__a21oi_2 _40905_ (.A1(_18309_),
    .A2(_18315_),
    .B1(_18316_),
    .Y(_18317_));
 sky130_fd_sc_hd__o211a_1 _40906_ (.A1(_18180_),
    .A2(_18195_),
    .B1(_18315_),
    .C1(_18309_),
    .X(_18318_));
 sky130_fd_sc_hd__o22ai_4 _40907_ (.A1(_18229_),
    .A2(_18230_),
    .B1(_18317_),
    .B2(_18318_),
    .Y(_18319_));
 sky130_fd_sc_hd__a21oi_1 _40908_ (.A1(_18312_),
    .A2(_18314_),
    .B1(_18313_),
    .Y(_18320_));
 sky130_fd_sc_hd__nor3_4 _40909_ (.A(_18308_),
    .B(_18299_),
    .C(_18300_),
    .Y(_18321_));
 sky130_fd_sc_hd__o21bai_2 _40910_ (.A1(_18320_),
    .A2(_18321_),
    .B1_N(_18316_),
    .Y(_18322_));
 sky130_fd_sc_hd__nand3_4 _40911_ (.A(_18309_),
    .B(_18316_),
    .C(_18315_),
    .Y(_18323_));
 sky130_fd_sc_hd__nor2_2 _40912_ (.A(_18230_),
    .B(_18229_),
    .Y(_18324_));
 sky130_fd_sc_hd__nand3_4 _40913_ (.A(_18322_),
    .B(_18323_),
    .C(_18324_),
    .Y(_18325_));
 sky130_fd_sc_hd__nand2_1 _40914_ (.A(_18192_),
    .B(_18211_),
    .Y(_18326_));
 sky130_fd_sc_hd__nand2_2 _40915_ (.A(_18326_),
    .B(_18197_),
    .Y(_18327_));
 sky130_fd_sc_hd__a21oi_4 _40916_ (.A1(_18319_),
    .A2(_18325_),
    .B1(_18327_),
    .Y(_18328_));
 sky130_fd_sc_hd__and3_1 _40917_ (.A(_18193_),
    .B(_18196_),
    .C(_18189_),
    .X(_18329_));
 sky130_fd_sc_hd__a31oi_1 _40918_ (.A1(_18188_),
    .A2(_18191_),
    .A3(_18190_),
    .B1(_18204_),
    .Y(_18330_));
 sky130_fd_sc_hd__o211a_2 _40919_ (.A1(_18329_),
    .A2(_18330_),
    .B1(_18325_),
    .C1(_18319_),
    .X(_18331_));
 sky130_fd_sc_hd__o22ai_4 _40920_ (.A1(_16818_),
    .A2(_18200_),
    .B1(_18328_),
    .B2(_18331_),
    .Y(_18332_));
 sky130_fd_sc_hd__a21oi_1 _40921_ (.A1(_18322_),
    .A2(_18323_),
    .B1(_18324_),
    .Y(_18333_));
 sky130_fd_sc_hd__nor2_1 _40922_ (.A(_17633_),
    .B(_18228_),
    .Y(_18334_));
 sky130_fd_sc_hd__nor2_1 _40923_ (.A(_16818_),
    .B(_18227_),
    .Y(_18335_));
 sky130_fd_sc_hd__o211a_1 _40924_ (.A1(_18334_),
    .A2(_18335_),
    .B1(_18323_),
    .C1(_18322_),
    .X(_18336_));
 sky130_fd_sc_hd__o21bai_2 _40925_ (.A1(_18333_),
    .A2(_18336_),
    .B1_N(_18327_),
    .Y(_18337_));
 sky130_fd_sc_hd__nand3_4 _40926_ (.A(_18319_),
    .B(_18327_),
    .C(_18325_),
    .Y(_18338_));
 sky130_fd_sc_hd__nand3_4 _40927_ (.A(_18337_),
    .B(_18207_),
    .C(_18338_),
    .Y(_18339_));
 sky130_vsdinv _40928_ (.A(_18094_),
    .Y(_18340_));
 sky130_fd_sc_hd__a21oi_2 _40929_ (.A1(_18210_),
    .A2(_18212_),
    .B1(_18120_),
    .Y(_18341_));
 sky130_fd_sc_hd__o21ai_4 _40930_ (.A1(_18340_),
    .A2(_18341_),
    .B1(_18213_),
    .Y(_18342_));
 sky130_fd_sc_hd__a21o_1 _40931_ (.A1(_18332_),
    .A2(_18339_),
    .B1(_18342_),
    .X(_18343_));
 sky130_fd_sc_hd__nand3_4 _40932_ (.A(_18332_),
    .B(_18342_),
    .C(_18339_),
    .Y(_18344_));
 sky130_fd_sc_hd__nand2_2 _40933_ (.A(_18343_),
    .B(_18344_),
    .Y(_18345_));
 sky130_vsdinv _40934_ (.A(_18219_),
    .Y(_18346_));
 sky130_fd_sc_hd__a21oi_4 _40935_ (.A1(_18226_),
    .A2(_18217_),
    .B1(_18346_),
    .Y(_18347_));
 sky130_fd_sc_hd__xor2_4 _40936_ (.A(_18345_),
    .B(_18347_),
    .X(_02680_));
 sky130_fd_sc_hd__nand2_2 _40937_ (.A(_18339_),
    .B(_18338_),
    .Y(_18348_));
 sky130_fd_sc_hd__a21oi_4 _40938_ (.A1(_18263_),
    .A2(_18255_),
    .B1(_18253_),
    .Y(_18349_));
 sky130_vsdinv _40939_ (.A(_18249_),
    .Y(_18350_));
 sky130_fd_sc_hd__nand2_4 _40940_ (.A(_18688_),
    .B(_16107_),
    .Y(_18351_));
 sky130_fd_sc_hd__or4_4 _40941_ (.A(_11607_),
    .B(_15914_),
    .C(_15916_),
    .D(_16147_),
    .X(_18352_));
 sky130_fd_sc_hd__a22o_1 _40942_ (.A1(_19831_),
    .A2(_10779_),
    .B1(_16059_),
    .B2(_15908_),
    .X(_18353_));
 sky130_fd_sc_hd__nand2_1 _40943_ (.A(_18352_),
    .B(_18353_),
    .Y(_18354_));
 sky130_fd_sc_hd__or2_2 _40944_ (.A(_18351_),
    .B(_18354_),
    .X(_18355_));
 sky130_fd_sc_hd__nand2_1 _40945_ (.A(_18354_),
    .B(_18351_),
    .Y(_18356_));
 sky130_fd_sc_hd__nand2_1 _40946_ (.A(_18355_),
    .B(_18356_),
    .Y(_18357_));
 sky130_fd_sc_hd__a21o_1 _40947_ (.A1(_18233_),
    .A2(_18236_),
    .B1(_18357_),
    .X(_18358_));
 sky130_fd_sc_hd__nand3_1 _40948_ (.A(_18357_),
    .B(_18233_),
    .C(_18236_),
    .Y(_18359_));
 sky130_fd_sc_hd__nand2_2 _40949_ (.A(_18358_),
    .B(_18359_),
    .Y(_18360_));
 sky130_fd_sc_hd__or2_4 _40950_ (.A(_18350_),
    .B(_18360_),
    .X(_18361_));
 sky130_fd_sc_hd__nand2_2 _40951_ (.A(_18360_),
    .B(_18350_),
    .Y(_18362_));
 sky130_fd_sc_hd__nor2_2 _40952_ (.A(_18238_),
    .B(_18242_),
    .Y(_18363_));
 sky130_fd_sc_hd__a21oi_4 _40953_ (.A1(_18243_),
    .A2(_18350_),
    .B1(_18363_),
    .Y(_18364_));
 sky130_fd_sc_hd__a21oi_4 _40954_ (.A1(_18361_),
    .A2(_18362_),
    .B1(_18364_),
    .Y(_18365_));
 sky130_fd_sc_hd__nand3_4 _40955_ (.A(_18361_),
    .B(_18364_),
    .C(_18362_),
    .Y(_18366_));
 sky130_vsdinv _40956_ (.A(_18366_),
    .Y(_18367_));
 sky130_vsdinv _40957_ (.A(_18033_),
    .Y(_18368_));
 sky130_vsdinv _40958_ (.A(_18245_),
    .Y(_18369_));
 sky130_fd_sc_hd__nand2_2 _40959_ (.A(_18247_),
    .B(_18369_),
    .Y(_18370_));
 sky130_vsdinv _40960_ (.A(_18370_),
    .Y(_18371_));
 sky130_fd_sc_hd__nand2_1 _40961_ (.A(_18368_),
    .B(_18371_),
    .Y(_18372_));
 sky130_fd_sc_hd__nand2_1 _40962_ (.A(_18033_),
    .B(_18370_),
    .Y(_18373_));
 sky130_fd_sc_hd__nand2_1 _40963_ (.A(_18372_),
    .B(_18373_),
    .Y(_18374_));
 sky130_fd_sc_hd__nor2_2 _40964_ (.A(_18030_),
    .B(_18374_),
    .Y(_18375_));
 sky130_fd_sc_hd__and2_1 _40965_ (.A(_18374_),
    .B(_18029_),
    .X(_18376_));
 sky130_fd_sc_hd__nor2_4 _40966_ (.A(_18375_),
    .B(_18376_),
    .Y(_18377_));
 sky130_vsdinv _40967_ (.A(_18377_),
    .Y(_18378_));
 sky130_fd_sc_hd__o21ai_2 _40968_ (.A1(_18365_),
    .A2(_18367_),
    .B1(_18378_),
    .Y(_18379_));
 sky130_fd_sc_hd__a21o_1 _40969_ (.A1(_18361_),
    .A2(_18362_),
    .B1(_18364_),
    .X(_18380_));
 sky130_fd_sc_hd__nand3_4 _40970_ (.A(_18380_),
    .B(_18366_),
    .C(_18377_),
    .Y(_18381_));
 sky130_fd_sc_hd__nand3b_4 _40971_ (.A_N(_18349_),
    .B(_18379_),
    .C(_18381_),
    .Y(_18382_));
 sky130_fd_sc_hd__o21ai_2 _40972_ (.A1(_18365_),
    .A2(_18367_),
    .B1(_18377_),
    .Y(_18383_));
 sky130_fd_sc_hd__nand3_2 _40973_ (.A(_18380_),
    .B(_18366_),
    .C(_18378_),
    .Y(_18384_));
 sky130_fd_sc_hd__nand3_4 _40974_ (.A(_18383_),
    .B(_18349_),
    .C(_18384_),
    .Y(_18385_));
 sky130_fd_sc_hd__nand2_2 _40975_ (.A(_18260_),
    .B(_18258_),
    .Y(_18386_));
 sky130_fd_sc_hd__xor2_4 _40976_ (.A(_17739_),
    .B(_18386_),
    .X(_18387_));
 sky130_fd_sc_hd__a21oi_2 _40977_ (.A1(_18382_),
    .A2(_18385_),
    .B1(_18387_),
    .Y(_18388_));
 sky130_fd_sc_hd__and3_1 _40978_ (.A(_18382_),
    .B(_18385_),
    .C(_18387_),
    .X(_18389_));
 sky130_fd_sc_hd__a21boi_2 _40979_ (.A1(_18270_),
    .A2(_18277_),
    .B1_N(_18267_),
    .Y(_18390_));
 sky130_fd_sc_hd__o21ai_4 _40980_ (.A1(_18388_),
    .A2(_18389_),
    .B1(_18390_),
    .Y(_18391_));
 sky130_fd_sc_hd__a21o_1 _40981_ (.A1(_18382_),
    .A2(_18385_),
    .B1(_18387_),
    .X(_18392_));
 sky130_fd_sc_hd__nand2_1 _40982_ (.A(_18280_),
    .B(_18267_),
    .Y(_18393_));
 sky130_fd_sc_hd__nand3_4 _40983_ (.A(_18382_),
    .B(_18385_),
    .C(_18387_),
    .Y(_18394_));
 sky130_fd_sc_hd__nand3_4 _40984_ (.A(_18392_),
    .B(_18393_),
    .C(_18394_),
    .Y(_18395_));
 sky130_fd_sc_hd__o21ai_2 _40985_ (.A1(_17844_),
    .A2(_18272_),
    .B1(_18274_),
    .Y(_18396_));
 sky130_vsdinv _40986_ (.A(_18396_),
    .Y(_18397_));
 sky130_fd_sc_hd__nand2_1 _40987_ (.A(_18397_),
    .B(_17315_),
    .Y(_18398_));
 sky130_fd_sc_hd__nand2_1 _40988_ (.A(_18396_),
    .B(_17316_),
    .Y(_18399_));
 sky130_fd_sc_hd__nand2_1 _40989_ (.A(_18398_),
    .B(_18399_),
    .Y(_18400_));
 sky130_fd_sc_hd__nand2_1 _40990_ (.A(_18397_),
    .B(_17314_),
    .Y(_18401_));
 sky130_fd_sc_hd__a21boi_4 _40991_ (.A1(_18401_),
    .A2(_16389_),
    .B1_N(_18399_),
    .Y(_18402_));
 sky130_fd_sc_hd__a22o_2 _40992_ (.A1(_17317_),
    .A2(_18400_),
    .B1(_18402_),
    .B2(_18398_),
    .X(_18403_));
 sky130_fd_sc_hd__a21oi_4 _40993_ (.A1(_18391_),
    .A2(_18395_),
    .B1(_18403_),
    .Y(_18404_));
 sky130_fd_sc_hd__and3_2 _40994_ (.A(_18391_),
    .B(_18395_),
    .C(_18403_),
    .X(_18405_));
 sky130_fd_sc_hd__a21boi_4 _40995_ (.A1(_18287_),
    .A2(_18295_),
    .B1_N(_18281_),
    .Y(_18406_));
 sky130_fd_sc_hd__o21ai_4 _40996_ (.A1(_18404_),
    .A2(_18405_),
    .B1(_18406_),
    .Y(_18407_));
 sky130_fd_sc_hd__nand2_2 _40997_ (.A(_18296_),
    .B(_18281_),
    .Y(_18408_));
 sky130_fd_sc_hd__a21o_1 _40998_ (.A1(_18391_),
    .A2(_18395_),
    .B1(_18403_),
    .X(_18409_));
 sky130_fd_sc_hd__nand3_4 _40999_ (.A(_18391_),
    .B(_18395_),
    .C(_18403_),
    .Y(_18410_));
 sky130_fd_sc_hd__nand3_4 _41000_ (.A(_18408_),
    .B(_18409_),
    .C(_18410_),
    .Y(_18411_));
 sky130_fd_sc_hd__nand2_1 _41001_ (.A(_18289_),
    .B(_17765_),
    .Y(_18412_));
 sky130_fd_sc_hd__nand2_1 _41002_ (.A(_18412_),
    .B(_18291_),
    .Y(_18413_));
 sky130_fd_sc_hd__or2_1 _41003_ (.A(_17944_),
    .B(_18413_),
    .X(_18414_));
 sky130_fd_sc_hd__nand2_1 _41004_ (.A(_18413_),
    .B(_17944_),
    .Y(_18415_));
 sky130_fd_sc_hd__a21oi_1 _41005_ (.A1(_18414_),
    .A2(_18415_),
    .B1(_17176_),
    .Y(_18416_));
 sky130_fd_sc_hd__and3_1 _41006_ (.A(_18414_),
    .B(_16992_),
    .C(_18415_),
    .X(_18417_));
 sky130_fd_sc_hd__or2_4 _41007_ (.A(_18416_),
    .B(_18417_),
    .X(_18418_));
 sky130_fd_sc_hd__a21oi_2 _41008_ (.A1(_18407_),
    .A2(_18411_),
    .B1(_18418_),
    .Y(_18419_));
 sky130_fd_sc_hd__and3_1 _41009_ (.A(_18407_),
    .B(_18418_),
    .C(_18411_),
    .X(_18420_));
 sky130_fd_sc_hd__o21ai_4 _41010_ (.A1(_18308_),
    .A2(_18299_),
    .B1(_18314_),
    .Y(_18421_));
 sky130_fd_sc_hd__o21bai_4 _41011_ (.A1(_18419_),
    .A2(_18420_),
    .B1_N(_18421_),
    .Y(_18422_));
 sky130_fd_sc_hd__a21oi_2 _41012_ (.A1(_18409_),
    .A2(_18410_),
    .B1(_18408_),
    .Y(_18423_));
 sky130_fd_sc_hd__nor3_4 _41013_ (.A(_18404_),
    .B(_18406_),
    .C(_18405_),
    .Y(_18424_));
 sky130_fd_sc_hd__o21bai_4 _41014_ (.A1(_18423_),
    .A2(_18424_),
    .B1_N(_18418_),
    .Y(_18425_));
 sky130_fd_sc_hd__nand3_4 _41015_ (.A(_18407_),
    .B(_18418_),
    .C(_18411_),
    .Y(_18426_));
 sky130_fd_sc_hd__nand3_4 _41016_ (.A(_18425_),
    .B(_18421_),
    .C(_18426_),
    .Y(_18427_));
 sky130_fd_sc_hd__and2_2 _41017_ (.A(_18305_),
    .B(_18302_),
    .X(_18428_));
 sky130_fd_sc_hd__nand2_4 _41018_ (.A(_18428_),
    .B(_17004_),
    .Y(_18429_));
 sky130_fd_sc_hd__a21o_1 _41019_ (.A1(_18305_),
    .A2(_18302_),
    .B1(_17004_),
    .X(_18430_));
 sky130_fd_sc_hd__and2_2 _41020_ (.A(_18429_),
    .B(_18430_),
    .X(_18431_));
 sky130_fd_sc_hd__a21bo_1 _41021_ (.A1(_18422_),
    .A2(_18427_),
    .B1_N(_18431_),
    .X(_18432_));
 sky130_fd_sc_hd__a31oi_4 _41022_ (.A1(_18425_),
    .A2(_18421_),
    .A3(_18426_),
    .B1(_18431_),
    .Y(_18433_));
 sky130_fd_sc_hd__nand2_2 _41023_ (.A(_18433_),
    .B(_18422_),
    .Y(_18434_));
 sky130_fd_sc_hd__nand2_2 _41024_ (.A(_18325_),
    .B(_18323_),
    .Y(_18435_));
 sky130_fd_sc_hd__a21oi_4 _41025_ (.A1(_18432_),
    .A2(_18434_),
    .B1(_18435_),
    .Y(_18436_));
 sky130_fd_sc_hd__and2_1 _41026_ (.A(_18325_),
    .B(_18323_),
    .X(_18437_));
 sky130_fd_sc_hd__nand2_1 _41027_ (.A(_18432_),
    .B(_18434_),
    .Y(_18438_));
 sky130_fd_sc_hd__nor2_1 _41028_ (.A(_18437_),
    .B(_18438_),
    .Y(_18439_));
 sky130_fd_sc_hd__or3_4 _41029_ (.A(_18229_),
    .B(_18436_),
    .C(_18439_),
    .X(_18440_));
 sky130_fd_sc_hd__or2_1 _41030_ (.A(_18437_),
    .B(_18438_),
    .X(_18441_));
 sky130_vsdinv _41031_ (.A(_18436_),
    .Y(_18442_));
 sky130_fd_sc_hd__nand2_1 _41032_ (.A(_18441_),
    .B(_18442_),
    .Y(_18443_));
 sky130_fd_sc_hd__nand2_1 _41033_ (.A(_18443_),
    .B(_18229_),
    .Y(_18444_));
 sky130_fd_sc_hd__nand3b_4 _41034_ (.A_N(_18348_),
    .B(_18440_),
    .C(_18444_),
    .Y(_18445_));
 sky130_vsdinv _41035_ (.A(_18229_),
    .Y(_18446_));
 sky130_fd_sc_hd__nand2_1 _41036_ (.A(_18443_),
    .B(_18446_),
    .Y(_18447_));
 sky130_fd_sc_hd__a21oi_2 _41037_ (.A1(_18438_),
    .A2(_18437_),
    .B1(_18446_),
    .Y(_18448_));
 sky130_fd_sc_hd__nand2_1 _41038_ (.A(_18441_),
    .B(_18448_),
    .Y(_18449_));
 sky130_fd_sc_hd__nand3_4 _41039_ (.A(_18447_),
    .B(_18348_),
    .C(_18449_),
    .Y(_18450_));
 sky130_fd_sc_hd__a21boi_4 _41040_ (.A1(_18219_),
    .A2(_18344_),
    .B1_N(_18343_),
    .Y(_18451_));
 sky130_vsdinv _41041_ (.A(_18207_),
    .Y(_18452_));
 sky130_fd_sc_hd__nor3_4 _41042_ (.A(_18452_),
    .B(_18328_),
    .C(_18331_),
    .Y(_18453_));
 sky130_fd_sc_hd__nand2_1 _41043_ (.A(_18332_),
    .B(_18342_),
    .Y(_18454_));
 sky130_fd_sc_hd__o2111ai_4 _41044_ (.A1(_18453_),
    .A2(_18454_),
    .B1(_18217_),
    .C1(_18219_),
    .D1(_18343_),
    .Y(_18455_));
 sky130_fd_sc_hd__a21oi_4 _41045_ (.A1(_18223_),
    .A2(_18225_),
    .B1(_18455_),
    .Y(_18456_));
 sky130_fd_sc_hd__a211oi_4 _41046_ (.A1(_18445_),
    .A2(_18450_),
    .B1(_18451_),
    .C1(_18456_),
    .Y(_18457_));
 sky130_fd_sc_hd__nand2_1 _41047_ (.A(_18445_),
    .B(_18450_),
    .Y(_18458_));
 sky130_fd_sc_hd__o21bai_2 _41048_ (.A1(_18451_),
    .A2(_18456_),
    .B1_N(_18458_),
    .Y(_18459_));
 sky130_fd_sc_hd__nor2b_1 _41049_ (.A(_18457_),
    .B_N(_18459_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor2_4 _41050_ (.A(_20071_),
    .B(_11276_),
    .Y(_18460_));
 sky130_fd_sc_hd__nand2_1 _41051_ (.A(_18410_),
    .B(_18395_),
    .Y(_18461_));
 sky130_fd_sc_hd__or2_2 _41052_ (.A(_18460_),
    .B(_18461_),
    .X(_18462_));
 sky130_fd_sc_hd__nand2_2 _41053_ (.A(_18461_),
    .B(_18460_),
    .Y(_18463_));
 sky130_fd_sc_hd__nand2_1 _41054_ (.A(_18381_),
    .B(_18380_),
    .Y(_18464_));
 sky130_vsdinv _41055_ (.A(_18464_),
    .Y(_18465_));
 sky130_fd_sc_hd__o21ai_4 _41056_ (.A1(_18249_),
    .A2(_18360_),
    .B1(_18358_),
    .Y(_18466_));
 sky130_fd_sc_hd__xnor2_2 _41057_ (.A(_18466_),
    .B(_18402_),
    .Y(_18467_));
 sky130_fd_sc_hd__xor2_4 _41058_ (.A(_18465_),
    .B(_18467_),
    .X(_18468_));
 sky130_fd_sc_hd__a21o_1 _41059_ (.A1(_18462_),
    .A2(_18463_),
    .B1(_18468_),
    .X(_18469_));
 sky130_fd_sc_hd__nand3_4 _41060_ (.A(_18462_),
    .B(_18468_),
    .C(_18463_),
    .Y(_18470_));
 sky130_fd_sc_hd__nand2_4 _41061_ (.A(_18355_),
    .B(_18352_),
    .Y(_18471_));
 sky130_fd_sc_hd__a21bo_2 _41062_ (.A1(_18414_),
    .A2(_17796_),
    .B1_N(_18415_),
    .X(_18472_));
 sky130_fd_sc_hd__xor2_4 _41063_ (.A(_18471_),
    .B(_18472_),
    .X(_18473_));
 sky130_fd_sc_hd__and3_1 _41064_ (.A(_18469_),
    .B(_18470_),
    .C(_18473_),
    .X(_18474_));
 sky130_fd_sc_hd__a21oi_4 _41065_ (.A1(_18469_),
    .A2(_18470_),
    .B1(_18473_),
    .Y(_18475_));
 sky130_fd_sc_hd__a31o_1 _41066_ (.A1(_18260_),
    .A2(_17737_),
    .A3(_18258_),
    .B1(_17735_),
    .X(_18476_));
 sky130_fd_sc_hd__xor2_4 _41067_ (.A(_18350_),
    .B(_18476_),
    .X(_18477_));
 sky130_fd_sc_hd__a21oi_4 _41068_ (.A1(_18425_),
    .A2(_18426_),
    .B1(_18421_),
    .Y(_18478_));
 sky130_fd_sc_hd__nor2_4 _41069_ (.A(_18429_),
    .B(_18478_),
    .Y(_18479_));
 sky130_fd_sc_hd__nand2_1 _41070_ (.A(_18427_),
    .B(_18429_),
    .Y(_18480_));
 sky130_fd_sc_hd__a21oi_4 _41071_ (.A1(_18433_),
    .A2(_18422_),
    .B1(_18480_),
    .Y(_18481_));
 sky130_fd_sc_hd__nor3_4 _41072_ (.A(_18477_),
    .B(_18479_),
    .C(_18481_),
    .Y(_18482_));
 sky130_fd_sc_hd__o211ai_4 _41073_ (.A1(_18431_),
    .A2(_18478_),
    .B1(_18427_),
    .C1(_18429_),
    .Y(_18483_));
 sky130_fd_sc_hd__nand3_4 _41074_ (.A(_18422_),
    .B(_17633_),
    .C(_18428_),
    .Y(_18484_));
 sky130_vsdinv _41075_ (.A(_18477_),
    .Y(_18485_));
 sky130_fd_sc_hd__a21oi_2 _41076_ (.A1(_18483_),
    .A2(_18484_),
    .B1(_18485_),
    .Y(_18486_));
 sky130_fd_sc_hd__o22ai_4 _41077_ (.A1(_18474_),
    .A2(_18475_),
    .B1(_18482_),
    .B2(_18486_),
    .Y(_18487_));
 sky130_fd_sc_hd__o21ai_2 _41078_ (.A1(_18479_),
    .A2(_18481_),
    .B1(_18477_),
    .Y(_18488_));
 sky130_fd_sc_hd__nor2_2 _41079_ (.A(_18475_),
    .B(_18474_),
    .Y(_18489_));
 sky130_fd_sc_hd__nand3_2 _41080_ (.A(_18483_),
    .B(_18485_),
    .C(_18484_),
    .Y(_18490_));
 sky130_fd_sc_hd__nand3_4 _41081_ (.A(_18488_),
    .B(_18489_),
    .C(_18490_),
    .Y(_18491_));
 sky130_vsdinv _41082_ (.A(_18434_),
    .Y(_18492_));
 sky130_fd_sc_hd__nand2_1 _41083_ (.A(_18432_),
    .B(_18435_),
    .Y(_18493_));
 sky130_fd_sc_hd__o22ai_4 _41084_ (.A1(_18492_),
    .A2(_18493_),
    .B1(_18446_),
    .B2(_18436_),
    .Y(_18494_));
 sky130_fd_sc_hd__a21oi_1 _41085_ (.A1(_18487_),
    .A2(_18491_),
    .B1(_18494_),
    .Y(_18495_));
 sky130_fd_sc_hd__o211a_1 _41086_ (.A1(_18439_),
    .A2(_18448_),
    .B1(_18491_),
    .C1(_18487_),
    .X(_18496_));
 sky130_fd_sc_hd__nand2_1 _41087_ (.A(_18394_),
    .B(_18382_),
    .Y(_18497_));
 sky130_fd_sc_hd__nand2_1 _41088_ (.A(_18426_),
    .B(_18411_),
    .Y(_18498_));
 sky130_fd_sc_hd__xor2_2 _41089_ (.A(_18351_),
    .B(_18498_),
    .X(_18499_));
 sky130_fd_sc_hd__xnor2_1 _41090_ (.A(_18497_),
    .B(_18499_),
    .Y(_18500_));
 sky130_fd_sc_hd__nor2_4 _41091_ (.A(_13024_),
    .B(_16103_),
    .Y(_18501_));
 sky130_fd_sc_hd__mux2_4 _41092_ (.A0(_16253_),
    .A1(_16252_),
    .S(_14014_),
    .X(_18502_));
 sky130_fd_sc_hd__xor2_4 _41093_ (.A(_18501_),
    .B(_18502_),
    .X(_18503_));
 sky130_fd_sc_hd__nand2_1 _41094_ (.A(_18500_),
    .B(_18503_),
    .Y(_18504_));
 sky130_fd_sc_hd__xor2_1 _41095_ (.A(_18497_),
    .B(_18499_),
    .X(_18505_));
 sky130_vsdinv _41096_ (.A(_18503_),
    .Y(_18506_));
 sky130_fd_sc_hd__nand2_1 _41097_ (.A(_18505_),
    .B(_18506_),
    .Y(_18507_));
 sky130_fd_sc_hd__nand2_1 _41098_ (.A(_18504_),
    .B(_18507_),
    .Y(_18508_));
 sky130_fd_sc_hd__o21bai_1 _41099_ (.A1(_18495_),
    .A2(_18496_),
    .B1_N(_18508_),
    .Y(_18509_));
 sky130_fd_sc_hd__a21o_1 _41100_ (.A1(_18487_),
    .A2(_18491_),
    .B1(_18494_),
    .X(_18510_));
 sky130_fd_sc_hd__nand3_1 _41101_ (.A(_18487_),
    .B(_18494_),
    .C(_18491_),
    .Y(_18511_));
 sky130_fd_sc_hd__nand3_2 _41102_ (.A(_18510_),
    .B(_18508_),
    .C(_18511_),
    .Y(_18512_));
 sky130_fd_sc_hd__nor2_2 _41103_ (.A(_18030_),
    .B(_18373_),
    .Y(_18513_));
 sky130_fd_sc_hd__and3_1 _41104_ (.A(_18368_),
    .B(_18030_),
    .C(_18371_),
    .X(_18514_));
 sky130_fd_sc_hd__or2_1 _41105_ (.A(_18513_),
    .B(_18514_),
    .X(_18515_));
 sky130_fd_sc_hd__a21oi_1 _41106_ (.A1(_18509_),
    .A2(_18512_),
    .B1(_18515_),
    .Y(_18516_));
 sky130_fd_sc_hd__o211a_1 _41107_ (.A1(_18513_),
    .A2(_18514_),
    .B1(_18512_),
    .C1(_18509_),
    .X(_18517_));
 sky130_fd_sc_hd__o2bb2ai_1 _41108_ (.A1_N(_18450_),
    .A2_N(_18459_),
    .B1(_18516_),
    .B2(_18517_),
    .Y(_18518_));
 sky130_fd_sc_hd__nor2_1 _41109_ (.A(_18516_),
    .B(_18517_),
    .Y(_18519_));
 sky130_fd_sc_hd__nand3_1 _41110_ (.A(_18519_),
    .B(_18450_),
    .C(_18459_),
    .Y(_18520_));
 sky130_fd_sc_hd__nand2_1 _41111_ (.A(_18518_),
    .B(_18520_),
    .Y(_02682_));
 sky130_fd_sc_hd__xor2_1 _41112_ (.A(_05358_),
    .B(_05210_),
    .X(_02628_));
 sky130_fd_sc_hd__nor2_1 _41113_ (.A(_20323_),
    .B(_04847_),
    .Y(_00050_));
 sky130_fd_sc_hd__and3_1 _41114_ (.A(_02321_),
    .B(_02318_),
    .C(_00066_),
    .X(_00068_));
 sky130_fd_sc_hd__and2_1 _41115_ (.A(_02321_),
    .B(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__and2_1 _41116_ (.A(_02321_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__o21a_4 _41117_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(net330),
    .X(_00216_));
 sky130_fd_sc_hd__o21a_1 _41118_ (.A1(_18748_),
    .A2(_18961_),
    .B1(_00321_),
    .X(_18521_));
 sky130_fd_sc_hd__nand2_1 _41119_ (.A(_18521_),
    .B(_18704_),
    .Y(_18522_));
 sky130_fd_sc_hd__o211a_1 _41120_ (.A1(irq_active),
    .A2(_18521_),
    .B1(_19195_),
    .C1(_18522_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _41121_ (.LO(net134));
 sky130_fd_sc_hd__conb_1 _41122_ (.LO(net145));
 sky130_fd_sc_hd__conb_1 _41123_ (.LO(net167));
 sky130_fd_sc_hd__conb_1 _41124_ (.LO(net178));
 sky130_fd_sc_hd__conb_1 _41125_ (.LO(net371));
 sky130_fd_sc_hd__conb_1 _41126_ (.LO(net382));
 sky130_fd_sc_hd__conb_1 _41127_ (.LO(net393));
 sky130_fd_sc_hd__conb_1 _41128_ (.LO(net400));
 sky130_fd_sc_hd__conb_1 _41129_ (.LO(net401));
 sky130_fd_sc_hd__conb_1 _41130_ (.LO(net402));
 sky130_fd_sc_hd__conb_1 _41131_ (.LO(net403));
 sky130_fd_sc_hd__conb_1 _41132_ (.LO(net404));
 sky130_fd_sc_hd__conb_1 _41133_ (.LO(net405));
 sky130_fd_sc_hd__conb_1 _41134_ (.LO(net406));
 sky130_fd_sc_hd__conb_1 _41135_ (.LO(net372));
 sky130_fd_sc_hd__conb_1 _41136_ (.LO(net373));
 sky130_fd_sc_hd__conb_1 _41137_ (.LO(net374));
 sky130_fd_sc_hd__conb_1 _41138_ (.LO(net375));
 sky130_fd_sc_hd__conb_1 _41139_ (.LO(net376));
 sky130_fd_sc_hd__conb_1 _41140_ (.LO(net377));
 sky130_fd_sc_hd__conb_1 _41141_ (.LO(net378));
 sky130_fd_sc_hd__conb_1 _41142_ (.LO(net379));
 sky130_fd_sc_hd__conb_1 _41143_ (.LO(net380));
 sky130_fd_sc_hd__conb_1 _41144_ (.LO(net381));
 sky130_fd_sc_hd__conb_1 _41145_ (.LO(net383));
 sky130_fd_sc_hd__conb_1 _41146_ (.LO(net384));
 sky130_fd_sc_hd__conb_1 _41147_ (.LO(net385));
 sky130_fd_sc_hd__conb_1 _41148_ (.LO(net386));
 sky130_fd_sc_hd__conb_1 _41149_ (.LO(net387));
 sky130_fd_sc_hd__conb_1 _41150_ (.LO(net388));
 sky130_fd_sc_hd__conb_1 _41151_ (.LO(net389));
 sky130_fd_sc_hd__conb_1 _41152_ (.LO(net390));
 sky130_fd_sc_hd__conb_1 _41153_ (.LO(net391));
 sky130_fd_sc_hd__conb_1 _41154_ (.LO(net392));
 sky130_fd_sc_hd__conb_1 _41155_ (.LO(net394));
 sky130_fd_sc_hd__conb_1 _41156_ (.LO(net395));
 sky130_fd_sc_hd__conb_1 _41157_ (.LO(net396));
 sky130_fd_sc_hd__conb_1 _41158_ (.LO(net397));
 sky130_fd_sc_hd__conb_1 _41159_ (.LO(net398));
 sky130_fd_sc_hd__conb_1 _41160_ (.LO(net399));
 sky130_fd_sc_hd__conb_1 _41161_ (.LO(net407));
 sky130_fd_sc_hd__conb_1 _41162_ (.LO(_00313_));
 sky130_fd_sc_hd__clkbuf_4 _41163_ (.A(net200),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 _41164_ (.A(net211),
    .X(net349));
 sky130_fd_sc_hd__buf_6 _41165_ (.A(net222),
    .X(net360));
 sky130_fd_sc_hd__buf_2 _41166_ (.A(net225),
    .X(net363));
 sky130_fd_sc_hd__buf_2 _41167_ (.A(net512),
    .X(net364));
 sky130_fd_sc_hd__buf_2 _41168_ (.A(net227),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _41169_ (.A(net228),
    .X(net366));
 sky130_fd_sc_hd__buf_2 _41170_ (.A(net229),
    .X(net367));
 sky130_fd_sc_hd__mux2_8 _41171_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(net459),
    .X(_21107_));
 sky130_fd_sc_hd__mux2_2 _41172_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_8 _41173_ (.A0(_02184_),
    .A1(net328),
    .S(net476),
    .X(net189));
 sky130_fd_sc_hd__mux2_2 _41174_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_8 _41175_ (.A0(_02185_),
    .A1(net331),
    .S(net476),
    .X(net192));
 sky130_fd_sc_hd__mux2_1 _41176_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_8 _41177_ (.A0(_02186_),
    .A1(net332),
    .S(net477),
    .X(net193));
 sky130_fd_sc_hd__mux2_1 _41178_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_8 _41179_ (.A0(_02187_),
    .A1(net333),
    .S(net477),
    .X(net194));
 sky130_fd_sc_hd__mux2_2 _41180_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_8 _41181_ (.A0(_02188_),
    .A1(net334),
    .S(net476),
    .X(net195));
 sky130_fd_sc_hd__mux2_2 _41182_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_8 _41183_ (.A0(_02189_),
    .A1(net335),
    .S(net476),
    .X(net196));
 sky130_fd_sc_hd__mux2_2 _41184_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_8 _41185_ (.A0(_02190_),
    .A1(net336),
    .S(net474),
    .X(net197));
 sky130_fd_sc_hd__mux2_1 _41186_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_8 _41187_ (.A0(_02191_),
    .A1(net337),
    .S(net477),
    .X(net198));
 sky130_fd_sc_hd__mux2_2 _41188_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_8 _41189_ (.A0(_02192_),
    .A1(net307),
    .S(net476),
    .X(net168));
 sky130_fd_sc_hd__mux2_2 _41190_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_8 _41191_ (.A0(_02193_),
    .A1(net308),
    .S(net476),
    .X(net169));
 sky130_fd_sc_hd__mux2_1 _41192_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_8 _41193_ (.A0(_02194_),
    .A1(net309),
    .S(net477),
    .X(net170));
 sky130_fd_sc_hd__mux2_2 _41194_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_8 _41195_ (.A0(_02195_),
    .A1(net310),
    .S(net476),
    .X(net171));
 sky130_fd_sc_hd__mux2_1 _41196_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_8 _41197_ (.A0(_02196_),
    .A1(net311),
    .S(net475),
    .X(net172));
 sky130_fd_sc_hd__mux2_1 _41198_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_2 _41199_ (.A0(_02197_),
    .A1(net312),
    .S(net474),
    .X(net173));
 sky130_fd_sc_hd__mux2_1 _41200_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_8 _41201_ (.A0(_02198_),
    .A1(net313),
    .S(net475),
    .X(net174));
 sky130_fd_sc_hd__mux2_1 _41202_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_8 _41203_ (.A0(_02199_),
    .A1(net314),
    .S(net475),
    .X(net175));
 sky130_fd_sc_hd__mux2_1 _41204_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_8 _41205_ (.A0(_02200_),
    .A1(net315),
    .S(net474),
    .X(net176));
 sky130_fd_sc_hd__mux2_1 _41206_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_8 _41207_ (.A0(_02201_),
    .A1(net316),
    .S(net474),
    .X(net177));
 sky130_fd_sc_hd__mux2_2 _41208_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_8 _41209_ (.A0(_02202_),
    .A1(net318),
    .S(net474),
    .X(net179));
 sky130_fd_sc_hd__mux2_1 _41210_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_8 _41211_ (.A0(_02203_),
    .A1(net319),
    .S(net475),
    .X(net180));
 sky130_fd_sc_hd__mux2_2 _41212_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_8 _41213_ (.A0(_02204_),
    .A1(net320),
    .S(net475),
    .X(net181));
 sky130_fd_sc_hd__mux2_2 _41214_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_8 _41215_ (.A0(_02205_),
    .A1(net321),
    .S(net474),
    .X(net182));
 sky130_fd_sc_hd__mux2_2 _41216_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_8 _41217_ (.A0(_02206_),
    .A1(net322),
    .S(net474),
    .X(net183));
 sky130_fd_sc_hd__mux2_2 _41218_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_4 _41219_ (.A0(_02207_),
    .A1(net323),
    .S(net474),
    .X(net184));
 sky130_fd_sc_hd__mux2_1 _41220_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_8 _41221_ (.A0(_02208_),
    .A1(net324),
    .S(net475),
    .X(net185));
 sky130_fd_sc_hd__mux2_1 _41222_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_4 _41223_ (.A0(_02209_),
    .A1(net325),
    .S(_00301_),
    .X(net186));
 sky130_fd_sc_hd__mux2_2 _41224_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_8 _41225_ (.A0(_02210_),
    .A1(net326),
    .S(net475),
    .X(net187));
 sky130_fd_sc_hd__mux2_1 _41226_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_8 _41227_ (.A0(_02211_),
    .A1(net327),
    .S(_00301_),
    .X(net188));
 sky130_fd_sc_hd__mux2_1 _41228_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_8 _41229_ (.A0(_02212_),
    .A1(net329),
    .S(_00301_),
    .X(net190));
 sky130_fd_sc_hd__mux2_4 _41230_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_4 _41231_ (.A0(_02213_),
    .A1(net330),
    .S(net474),
    .X(net191));
 sky130_fd_sc_hd__mux2_8 _41232_ (.A0(_02167_),
    .A1(net368),
    .S(_01683_),
    .X(net230));
 sky130_fd_sc_hd__mux2_8 _41233_ (.A0(_02168_),
    .A1(net369),
    .S(net452),
    .X(net231));
 sky130_fd_sc_hd__mux2_8 _41234_ (.A0(_02169_),
    .A1(net339),
    .S(_01683_),
    .X(net201));
 sky130_fd_sc_hd__mux2_8 _41235_ (.A0(_02170_),
    .A1(net340),
    .S(net452),
    .X(net202));
 sky130_fd_sc_hd__mux2_8 _41236_ (.A0(_02171_),
    .A1(net341),
    .S(net451),
    .X(net203));
 sky130_fd_sc_hd__mux2_4 _41237_ (.A0(_02172_),
    .A1(net342),
    .S(net452),
    .X(net204));
 sky130_fd_sc_hd__mux2_8 _41238_ (.A0(_02173_),
    .A1(net343),
    .S(net451),
    .X(net205));
 sky130_fd_sc_hd__mux2_8 _41239_ (.A0(_02174_),
    .A1(net344),
    .S(net451),
    .X(net206));
 sky130_fd_sc_hd__mux2_8 _41240_ (.A0(_02175_),
    .A1(net345),
    .S(net450),
    .X(net207));
 sky130_fd_sc_hd__mux2_8 _41241_ (.A0(_02176_),
    .A1(net346),
    .S(net453),
    .X(net208));
 sky130_fd_sc_hd__mux2_8 _41242_ (.A0(_02177_),
    .A1(net347),
    .S(net452),
    .X(net209));
 sky130_fd_sc_hd__mux2_8 _41243_ (.A0(_02178_),
    .A1(net348),
    .S(net452),
    .X(net210));
 sky130_fd_sc_hd__mux2_8 _41244_ (.A0(_02179_),
    .A1(net350),
    .S(net452),
    .X(net212));
 sky130_fd_sc_hd__mux2_8 _41245_ (.A0(_02180_),
    .A1(net351),
    .S(net453),
    .X(net213));
 sky130_fd_sc_hd__mux2_8 _41246_ (.A0(_02181_),
    .A1(net352),
    .S(net453),
    .X(net214));
 sky130_fd_sc_hd__mux2_8 _41247_ (.A0(_02182_),
    .A1(net353),
    .S(net453),
    .X(net215));
 sky130_fd_sc_hd__mux2_8 _41248_ (.A0(_02167_),
    .A1(net354),
    .S(_01683_),
    .X(net216));
 sky130_fd_sc_hd__mux2_8 _41249_ (.A0(_02168_),
    .A1(net355),
    .S(net452),
    .X(net217));
 sky130_fd_sc_hd__mux2_8 _41250_ (.A0(_02169_),
    .A1(net356),
    .S(_01683_),
    .X(net218));
 sky130_fd_sc_hd__mux2_8 _41251_ (.A0(_02170_),
    .A1(net357),
    .S(net452),
    .X(net219));
 sky130_fd_sc_hd__mux2_4 _41252_ (.A0(_02171_),
    .A1(net358),
    .S(net451),
    .X(net220));
 sky130_fd_sc_hd__mux2_8 _41253_ (.A0(_02172_),
    .A1(net359),
    .S(net452),
    .X(net221));
 sky130_fd_sc_hd__mux2_8 _41254_ (.A0(_02173_),
    .A1(net361),
    .S(net451),
    .X(net223));
 sky130_fd_sc_hd__mux2_4 _41255_ (.A0(_02174_),
    .A1(net362),
    .S(net451),
    .X(net224));
 sky130_fd_sc_hd__mux2_1 _41256_ (.A0(\mem_rdata_q[7] ),
    .A1(net62),
    .S(mem_xfer),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _41257_ (.A0(\mem_rdata_q[8] ),
    .A1(net63),
    .S(net437),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _41258_ (.A0(\mem_rdata_q[9] ),
    .A1(net64),
    .S(net437),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _41259_ (.A0(\mem_rdata_q[10] ),
    .A1(net34),
    .S(net437),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _41260_ (.A0(\mem_rdata_q[11] ),
    .A1(net35),
    .S(net437),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_2 _41261_ (.A0(\mem_rdata_q[12] ),
    .A1(net528),
    .S(net437),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_2 _41262_ (.A0(\mem_rdata_q[13] ),
    .A1(net37),
    .S(net437),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_2 _41263_ (.A0(\mem_rdata_q[14] ),
    .A1(net38),
    .S(net437),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_1 _41264_ (.A0(\mem_rdata_q[15] ),
    .A1(net527),
    .S(net437),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _41265_ (.A0(\mem_rdata_q[16] ),
    .A1(net40),
    .S(net437),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _41266_ (.A0(\mem_rdata_q[17] ),
    .A1(net41),
    .S(net437),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _41267_ (.A0(\mem_rdata_q[18] ),
    .A1(net42),
    .S(net437),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _41268_ (.A0(\mem_rdata_q[19] ),
    .A1(net526),
    .S(net437),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _41269_ (.A0(\mem_rdata_q[20] ),
    .A1(net524),
    .S(net437),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _41270_ (.A0(\mem_rdata_q[21] ),
    .A1(net46),
    .S(net437),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _41271_ (.A0(\mem_rdata_q[22] ),
    .A1(net47),
    .S(net437),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _41272_ (.A0(\mem_rdata_q[23] ),
    .A1(net48),
    .S(mem_xfer),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _41273_ (.A0(\mem_rdata_q[24] ),
    .A1(net49),
    .S(net437),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_1 _41274_ (.A0(\mem_rdata_q[25] ),
    .A1(net50),
    .S(mem_xfer),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_1 _41275_ (.A0(\mem_rdata_q[26] ),
    .A1(net51),
    .S(net437),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_1 _41276_ (.A0(\mem_rdata_q[27] ),
    .A1(net52),
    .S(mem_xfer),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_1 _41277_ (.A0(\mem_rdata_q[28] ),
    .A1(net53),
    .S(mem_xfer),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _41278_ (.A0(\mem_rdata_q[29] ),
    .A1(net54),
    .S(net437),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _41279_ (.A0(\mem_rdata_q[30] ),
    .A1(net523),
    .S(net437),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_1 _41280_ (.A0(\mem_rdata_q[31] ),
    .A1(net57),
    .S(mem_xfer),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _41281_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _41282_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _41283_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _41284_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _41285_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _41286_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _41287_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _41288_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _41289_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _41290_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _41291_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _41292_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_1 _41293_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _41294_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _41295_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _41296_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _41297_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _41298_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _41299_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _41300_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_1 _41301_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _41302_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _41303_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_1 _41304_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_1 _41305_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_1 _41306_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_1 _41307_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _41308_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_1 _41309_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_1 _41310_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_1 _41311_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_1 _41312_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_4 _41313_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_8 _41314_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(net431),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_8 _41315_ (.A0(_02074_),
    .A1(_02073_),
    .S(net429),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_8 _41316_ (.A0(_02076_),
    .A1(_02075_),
    .S(net429),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_8 _41317_ (.A0(_02078_),
    .A1(_02077_),
    .S(net429),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_8 _41318_ (.A0(_02080_),
    .A1(_02079_),
    .S(net429),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_8 _41319_ (.A0(_02082_),
    .A1(_02081_),
    .S(net429),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_8 _41320_ (.A0(_02084_),
    .A1(_02083_),
    .S(net429),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_8 _41321_ (.A0(_02086_),
    .A1(_02085_),
    .S(net429),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_8 _41322_ (.A0(_02088_),
    .A1(_02087_),
    .S(net429),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_8 _41323_ (.A0(_02090_),
    .A1(_02089_),
    .S(net429),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_8 _41324_ (.A0(_02092_),
    .A1(_02091_),
    .S(net431),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_4 _41325_ (.A0(_02094_),
    .A1(_02093_),
    .S(net431),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_4 _41326_ (.A0(_02096_),
    .A1(_02095_),
    .S(net431),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_4 _41327_ (.A0(_02098_),
    .A1(_02097_),
    .S(net431),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_2 _41328_ (.A0(_02100_),
    .A1(_02099_),
    .S(net430),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_4 _41329_ (.A0(_02102_),
    .A1(_02101_),
    .S(net430),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_4 _41330_ (.A0(_02104_),
    .A1(_02103_),
    .S(net430),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_4 _41331_ (.A0(_02106_),
    .A1(_02105_),
    .S(net430),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_4 _41332_ (.A0(_02108_),
    .A1(_02107_),
    .S(net430),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_2 _41333_ (.A0(_02110_),
    .A1(_02109_),
    .S(net430),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_2 _41334_ (.A0(_02112_),
    .A1(_02111_),
    .S(net430),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_2 _41335_ (.A0(_02114_),
    .A1(_02113_),
    .S(net430),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_4 _41336_ (.A0(_02116_),
    .A1(_02115_),
    .S(net430),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_4 _41337_ (.A0(_02118_),
    .A1(_02117_),
    .S(net430),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_4 _41338_ (.A0(_02120_),
    .A1(_02119_),
    .S(net430),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_4 _41339_ (.A0(_02122_),
    .A1(_02121_),
    .S(net430),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_2 _41340_ (.A0(_02124_),
    .A1(_02123_),
    .S(net430),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_2 _41341_ (.A0(_02126_),
    .A1(_02125_),
    .S(net430),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_4 _41342_ (.A0(_02128_),
    .A1(_02127_),
    .S(net431),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_2 _41343_ (.A0(_02130_),
    .A1(_02129_),
    .S(net431),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_2 _41344_ (.A0(_02132_),
    .A1(_02131_),
    .S(net431),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _41345_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _41346_ (.A0(_00347_),
    .A1(_21108_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _41347_ (.A0(_21108_),
    .A1(_00348_),
    .S(net101),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _41348_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _41349_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _41350_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _41351_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _41352_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _41353_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _41354_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _41355_ (.A0(_02223_),
    .A1(_02221_),
    .S(_02217_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _41356_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _41357_ (.A0(_02226_),
    .A1(_02224_),
    .S(net428),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _41358_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _41359_ (.A0(_02229_),
    .A1(_02227_),
    .S(net428),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _41360_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _41361_ (.A0(_02232_),
    .A1(_02230_),
    .S(net428),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _41362_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _41363_ (.A0(_02235_),
    .A1(_02233_),
    .S(net428),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _41364_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _41365_ (.A0(_02238_),
    .A1(_02236_),
    .S(net428),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _41366_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _41367_ (.A0(_02241_),
    .A1(_02239_),
    .S(net428),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _41368_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _41369_ (.A0(_02244_),
    .A1(_02242_),
    .S(net428),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _41370_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _41371_ (.A0(_02247_),
    .A1(_02245_),
    .S(_02217_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _41372_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _41373_ (.A0(_02250_),
    .A1(_02248_),
    .S(net428),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _41374_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _41375_ (.A0(_02253_),
    .A1(_02251_),
    .S(net428),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _41376_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _41377_ (.A0(_02256_),
    .A1(_02254_),
    .S(net428),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _41378_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _41379_ (.A0(_02259_),
    .A1(_02257_),
    .S(net428),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _41380_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _41381_ (.A0(_02262_),
    .A1(_02260_),
    .S(net428),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _41382_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _41383_ (.A0(_02265_),
    .A1(_02263_),
    .S(net428),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _41384_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _41385_ (.A0(_02268_),
    .A1(_02266_),
    .S(net428),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _41386_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _41387_ (.A0(_02271_),
    .A1(_02269_),
    .S(net428),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _41388_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _41389_ (.A0(_02274_),
    .A1(_02272_),
    .S(net428),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _41390_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _41391_ (.A0(_02277_),
    .A1(_02275_),
    .S(net428),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _41392_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _41393_ (.A0(_02280_),
    .A1(_02278_),
    .S(net428),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _41394_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _41395_ (.A0(_02283_),
    .A1(_02281_),
    .S(net428),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _41396_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _41397_ (.A0(_02286_),
    .A1(_02284_),
    .S(net428),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _41398_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _41399_ (.A0(_02289_),
    .A1(_02287_),
    .S(net428),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _41400_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _41401_ (.A0(_02292_),
    .A1(_02290_),
    .S(net428),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _41402_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _41403_ (.A0(_02295_),
    .A1(_02293_),
    .S(net428),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _41404_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _41405_ (.A0(_02298_),
    .A1(_02296_),
    .S(net428),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _41406_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _41407_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_2 _41408_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(net472),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_2 _41409_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(net472),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_4 _41410_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(net472),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_2 _41411_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(net472),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_2 _41412_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(net472),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_2 _41413_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(net472),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_2 _41414_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(net472),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_4 _41415_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(net472),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_2 _41416_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(net472),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_2 _41417_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(net472),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_2 _41418_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(net472),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_2 _41419_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(net472),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_2 _41420_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(net472),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_2 _41421_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(net471),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_2 _41422_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(net471),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_2 _41423_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(net471),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_2 _41424_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(net471),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_2 _41425_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(net471),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_2 _41426_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(net471),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_2 _41427_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(net471),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_4 _41428_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(net471),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_2 _41429_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(net471),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_4 _41430_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(net471),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_4 _41431_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(net471),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_4 _41432_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(net471),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_2 _41433_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(net471),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_4 _41434_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(net471),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_2 _41435_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(net471),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_4 _41436_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(_00292_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_2 _41437_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _41438_ (.A0(_00057_),
    .A1(_00064_),
    .S(net225),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _41439_ (.A0(_00065_),
    .A1(_02543_),
    .S(net226),
    .X(_21144_));
 sky130_fd_sc_hd__mux2_1 _41440_ (.A0(_00075_),
    .A1(_00082_),
    .S(net513),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _41441_ (.A0(_00083_),
    .A1(_02544_),
    .S(net512),
    .X(_21145_));
 sky130_fd_sc_hd__mux2_1 _41442_ (.A0(_00089_),
    .A1(_00092_),
    .S(net225),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _41443_ (.A0(_00093_),
    .A1(_02545_),
    .S(net226),
    .X(_21146_));
 sky130_fd_sc_hd__mux2_1 _41444_ (.A0(_00099_),
    .A1(_00102_),
    .S(net513),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _41445_ (.A0(_00103_),
    .A1(_02546_),
    .S(net512),
    .X(_21147_));
 sky130_fd_sc_hd__mux2_1 _41446_ (.A0(_00107_),
    .A1(_00108_),
    .S(net225),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _41447_ (.A0(_00109_),
    .A1(_02547_),
    .S(net226),
    .X(_21148_));
 sky130_fd_sc_hd__mux2_1 _41448_ (.A0(_00113_),
    .A1(_00114_),
    .S(net513),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _41449_ (.A0(_00115_),
    .A1(_02548_),
    .S(net512),
    .X(_21149_));
 sky130_fd_sc_hd__mux2_1 _41450_ (.A0(_00119_),
    .A1(_00120_),
    .S(net225),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _41451_ (.A0(_00121_),
    .A1(_02549_),
    .S(net512),
    .X(_21150_));
 sky130_fd_sc_hd__mux2_1 _41452_ (.A0(_00125_),
    .A1(_00126_),
    .S(net513),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _41453_ (.A0(_00127_),
    .A1(_02550_),
    .S(net512),
    .X(_21151_));
 sky130_fd_sc_hd__mux2_1 _41454_ (.A0(_00129_),
    .A1(_00106_),
    .S(net222),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _41455_ (.A0(_00130_),
    .A1(_00057_),
    .S(net225),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _41456_ (.A0(_00131_),
    .A1(_02551_),
    .S(net226),
    .X(_21152_));
 sky130_fd_sc_hd__mux2_1 _41457_ (.A0(_00133_),
    .A1(_00112_),
    .S(net514),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _41458_ (.A0(_00134_),
    .A1(_00075_),
    .S(net513),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _41459_ (.A0(_00135_),
    .A1(_02552_),
    .S(net512),
    .X(_21153_));
 sky130_fd_sc_hd__mux2_1 _41460_ (.A0(_00137_),
    .A1(_00118_),
    .S(net222),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _41461_ (.A0(_00138_),
    .A1(_00089_),
    .S(net225),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _41462_ (.A0(_00139_),
    .A1(_02553_),
    .S(net512),
    .X(_21154_));
 sky130_fd_sc_hd__mux2_1 _41463_ (.A0(_00141_),
    .A1(_00124_),
    .S(net514),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _41464_ (.A0(_00142_),
    .A1(_00099_),
    .S(net513),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _41465_ (.A0(_00143_),
    .A1(_02554_),
    .S(net512),
    .X(_21155_));
 sky130_fd_sc_hd__mux2_1 _41466_ (.A0(_00144_),
    .A1(_00136_),
    .S(net211),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _41467_ (.A0(_00145_),
    .A1(_00129_),
    .S(net222),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _41468_ (.A0(_00146_),
    .A1(_00107_),
    .S(net225),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _41469_ (.A0(_00147_),
    .A1(_02555_),
    .S(net226),
    .X(_21156_));
 sky130_fd_sc_hd__mux2_1 _41470_ (.A0(_00148_),
    .A1(_00140_),
    .S(net515),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _41471_ (.A0(_00149_),
    .A1(_00133_),
    .S(net514),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _41472_ (.A0(_00150_),
    .A1(_00113_),
    .S(net513),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _41473_ (.A0(_00151_),
    .A1(_02556_),
    .S(net512),
    .X(_21157_));
 sky130_fd_sc_hd__mux2_1 _41474_ (.A0(net329),
    .A1(net327),
    .S(net200),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _41475_ (.A0(_00152_),
    .A1(_00144_),
    .S(net211),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _41476_ (.A0(_00153_),
    .A1(_00137_),
    .S(net222),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _41477_ (.A0(_00154_),
    .A1(_00119_),
    .S(net225),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _41478_ (.A0(_00155_),
    .A1(_02557_),
    .S(net512),
    .X(_21158_));
 sky130_fd_sc_hd__mux2_1 _41479_ (.A0(net330),
    .A1(net329),
    .S(net516),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _41480_ (.A0(_00156_),
    .A1(_00148_),
    .S(net515),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _41481_ (.A0(_00157_),
    .A1(_00141_),
    .S(net514),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _41482_ (.A0(_00158_),
    .A1(_00125_),
    .S(net513),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _41483_ (.A0(_00159_),
    .A1(_02558_),
    .S(net512),
    .X(_21159_));
 sky130_fd_sc_hd__mux2_1 _41484_ (.A0(net306),
    .A1(net317),
    .S(net516),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _41485_ (.A0(_00160_),
    .A1(_00161_),
    .S(net515),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _41486_ (.A0(_00162_),
    .A1(_00165_),
    .S(net514),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _41487_ (.A0(_00166_),
    .A1(_00173_),
    .S(net513),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_2 _41488_ (.A0(_00174_),
    .A1(_00189_),
    .S(net512),
    .X(_21160_));
 sky130_fd_sc_hd__mux2_1 _41489_ (.A0(net317),
    .A1(net328),
    .S(net516),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _41490_ (.A0(_00190_),
    .A1(_00191_),
    .S(net515),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _41491_ (.A0(_00192_),
    .A1(_00195_),
    .S(net514),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _41492_ (.A0(_00196_),
    .A1(_00203_),
    .S(net513),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _41493_ (.A0(_00204_),
    .A1(_00220_),
    .S(net512),
    .X(_21171_));
 sky130_fd_sc_hd__mux2_1 _41494_ (.A0(_00161_),
    .A1(_00163_),
    .S(net515),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _41495_ (.A0(_00221_),
    .A1(_00222_),
    .S(net514),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _41496_ (.A0(_00223_),
    .A1(_00226_),
    .S(net513),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _41497_ (.A0(_00227_),
    .A1(_00234_),
    .S(net512),
    .X(_21182_));
 sky130_fd_sc_hd__mux2_1 _41498_ (.A0(_00191_),
    .A1(_00193_),
    .S(net515),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _41499_ (.A0(_00235_),
    .A1(_00236_),
    .S(net514),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _41500_ (.A0(_00237_),
    .A1(_00240_),
    .S(net513),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _41501_ (.A0(_00241_),
    .A1(_00248_),
    .S(net512),
    .X(_21185_));
 sky130_fd_sc_hd__mux2_1 _41502_ (.A0(_00165_),
    .A1(_00169_),
    .S(net514),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _41503_ (.A0(_00249_),
    .A1(_00250_),
    .S(net513),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _41504_ (.A0(_00251_),
    .A1(_00254_),
    .S(net512),
    .X(_21186_));
 sky130_fd_sc_hd__mux2_1 _41505_ (.A0(_00195_),
    .A1(_00199_),
    .S(net514),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _41506_ (.A0(_00255_),
    .A1(_00256_),
    .S(net513),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _41507_ (.A0(_00257_),
    .A1(_00260_),
    .S(net512),
    .X(_21187_));
 sky130_fd_sc_hd__mux2_1 _41508_ (.A0(_00222_),
    .A1(_00224_),
    .S(net514),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _41509_ (.A0(_00261_),
    .A1(_00262_),
    .S(net513),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _41510_ (.A0(_00263_),
    .A1(_00266_),
    .S(net512),
    .X(_21188_));
 sky130_fd_sc_hd__mux2_1 _41511_ (.A0(_00236_),
    .A1(_00238_),
    .S(net514),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _41512_ (.A0(_00267_),
    .A1(_00268_),
    .S(net513),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _41513_ (.A0(_00269_),
    .A1(_00272_),
    .S(net512),
    .X(_21189_));
 sky130_fd_sc_hd__mux2_1 _41514_ (.A0(_00173_),
    .A1(_00181_),
    .S(net513),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _41515_ (.A0(_00273_),
    .A1(_00274_),
    .S(net512),
    .X(_21190_));
 sky130_fd_sc_hd__mux2_1 _41516_ (.A0(_00203_),
    .A1(_00211_),
    .S(net513),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _41517_ (.A0(_00275_),
    .A1(_00276_),
    .S(net512),
    .X(_21191_));
 sky130_fd_sc_hd__mux2_1 _41518_ (.A0(_00226_),
    .A1(_00230_),
    .S(net513),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _41519_ (.A0(_00277_),
    .A1(_00278_),
    .S(net512),
    .X(_21161_));
 sky130_fd_sc_hd__mux2_1 _41520_ (.A0(_00240_),
    .A1(_00244_),
    .S(net513),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _41521_ (.A0(_00279_),
    .A1(_00280_),
    .S(net512),
    .X(_21162_));
 sky130_fd_sc_hd__mux2_1 _41522_ (.A0(_00250_),
    .A1(_00252_),
    .S(net513),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _41523_ (.A0(_00281_),
    .A1(_00282_),
    .S(net512),
    .X(_21163_));
 sky130_fd_sc_hd__mux2_1 _41524_ (.A0(_00256_),
    .A1(_00258_),
    .S(net513),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _41525_ (.A0(_00283_),
    .A1(_00284_),
    .S(net512),
    .X(_21164_));
 sky130_fd_sc_hd__mux2_1 _41526_ (.A0(_00262_),
    .A1(_00264_),
    .S(net513),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _41527_ (.A0(_00285_),
    .A1(_00286_),
    .S(net512),
    .X(_21165_));
 sky130_fd_sc_hd__mux2_1 _41528_ (.A0(_00268_),
    .A1(_00270_),
    .S(net513),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _41529_ (.A0(_00287_),
    .A1(_00288_),
    .S(net512),
    .X(_21166_));
 sky130_fd_sc_hd__mux2_1 _41530_ (.A0(_00189_),
    .A1(_00216_),
    .S(net512),
    .X(_21167_));
 sky130_fd_sc_hd__mux2_1 _41531_ (.A0(_00220_),
    .A1(_00216_),
    .S(net512),
    .X(_21168_));
 sky130_fd_sc_hd__mux2_1 _41532_ (.A0(_00234_),
    .A1(_00216_),
    .S(net512),
    .X(_21169_));
 sky130_fd_sc_hd__mux2_1 _41533_ (.A0(_00248_),
    .A1(_00216_),
    .S(net512),
    .X(_21170_));
 sky130_fd_sc_hd__mux2_1 _41534_ (.A0(_00254_),
    .A1(_00216_),
    .S(net512),
    .X(_21172_));
 sky130_fd_sc_hd__mux2_1 _41535_ (.A0(_00260_),
    .A1(_00216_),
    .S(net512),
    .X(_21173_));
 sky130_fd_sc_hd__mux2_1 _41536_ (.A0(_00266_),
    .A1(_00216_),
    .S(net512),
    .X(_21174_));
 sky130_fd_sc_hd__mux2_1 _41537_ (.A0(_00272_),
    .A1(_00216_),
    .S(net512),
    .X(_21175_));
 sky130_fd_sc_hd__mux2_1 _41538_ (.A0(_00274_),
    .A1(_00216_),
    .S(net512),
    .X(_21176_));
 sky130_fd_sc_hd__mux2_1 _41539_ (.A0(_00276_),
    .A1(_00216_),
    .S(net512),
    .X(_21177_));
 sky130_fd_sc_hd__mux2_1 _41540_ (.A0(_00278_),
    .A1(_00216_),
    .S(net512),
    .X(_21178_));
 sky130_fd_sc_hd__mux2_1 _41541_ (.A0(_00280_),
    .A1(_00216_),
    .S(net512),
    .X(_21179_));
 sky130_fd_sc_hd__mux2_1 _41542_ (.A0(_00282_),
    .A1(_00216_),
    .S(net512),
    .X(_21180_));
 sky130_fd_sc_hd__mux2_1 _41543_ (.A0(_00284_),
    .A1(_00216_),
    .S(net512),
    .X(_21181_));
 sky130_fd_sc_hd__mux2_1 _41544_ (.A0(_00286_),
    .A1(_00216_),
    .S(net512),
    .X(_21183_));
 sky130_fd_sc_hd__mux2_1 _41545_ (.A0(_00288_),
    .A1(_00216_),
    .S(net512),
    .X(_21184_));
 sky130_fd_sc_hd__mux2_1 _41546_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _41547_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_21143_));
 sky130_fd_sc_hd__mux2_1 _41548_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_21109_));
 sky130_fd_sc_hd__mux2_1 _41549_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(_01706_),
    .X(_21120_));
 sky130_fd_sc_hd__mux2_1 _41550_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(_01706_),
    .X(_21131_));
 sky130_fd_sc_hd__mux2_1 _41551_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(_01706_),
    .X(_21134_));
 sky130_fd_sc_hd__mux2_1 _41552_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(_01706_),
    .X(_21135_));
 sky130_fd_sc_hd__mux2_1 _41553_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(_01706_),
    .X(_21136_));
 sky130_fd_sc_hd__mux2_1 _41554_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(_01706_),
    .X(_21137_));
 sky130_fd_sc_hd__mux2_1 _41555_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(_01706_),
    .X(_21138_));
 sky130_fd_sc_hd__mux2_1 _41556_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(_01706_),
    .X(_21139_));
 sky130_fd_sc_hd__mux2_1 _41557_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(_01706_),
    .X(_21140_));
 sky130_fd_sc_hd__mux2_1 _41558_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(_01706_),
    .X(_21110_));
 sky130_fd_sc_hd__mux2_1 _41559_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(_01706_),
    .X(_21111_));
 sky130_fd_sc_hd__mux2_1 _41560_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(_01706_),
    .X(_21112_));
 sky130_fd_sc_hd__mux2_1 _41561_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(_01706_),
    .X(_21113_));
 sky130_fd_sc_hd__mux2_1 _41562_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(_01706_),
    .X(_21114_));
 sky130_fd_sc_hd__mux2_2 _41563_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(_01706_),
    .X(_21115_));
 sky130_fd_sc_hd__mux2_1 _41564_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(_01706_),
    .X(_21116_));
 sky130_fd_sc_hd__mux2_1 _41565_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(_01706_),
    .X(_21117_));
 sky130_fd_sc_hd__mux2_1 _41566_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(_01706_),
    .X(_21118_));
 sky130_fd_sc_hd__mux2_1 _41567_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(_01706_),
    .X(_21119_));
 sky130_fd_sc_hd__mux2_1 _41568_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(_01706_),
    .X(_21121_));
 sky130_fd_sc_hd__mux2_1 _41569_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(_01706_),
    .X(_21122_));
 sky130_fd_sc_hd__mux2_1 _41570_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(_01706_),
    .X(_21123_));
 sky130_fd_sc_hd__mux2_1 _41571_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(_01706_),
    .X(_21124_));
 sky130_fd_sc_hd__mux2_1 _41572_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(_01706_),
    .X(_21125_));
 sky130_fd_sc_hd__mux2_1 _41573_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(_01706_),
    .X(_21126_));
 sky130_fd_sc_hd__mux2_1 _41574_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(_01706_),
    .X(_21127_));
 sky130_fd_sc_hd__mux2_1 _41575_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_21128_));
 sky130_fd_sc_hd__mux2_1 _41576_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(_01706_),
    .X(_21129_));
 sky130_fd_sc_hd__mux2_1 _41577_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_21130_));
 sky130_fd_sc_hd__mux2_1 _41578_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_21132_));
 sky130_fd_sc_hd__mux2_1 _41579_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(_01706_),
    .X(_21133_));
 sky130_fd_sc_hd__mux2_1 _41580_ (.A0(_02061_),
    .A1(net518),
    .S(_02542_),
    .X(_21104_));
 sky130_fd_sc_hd__mux2_8 _41581_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(_00308_),
    .X(_21103_));
 sky130_fd_sc_hd__mux2_1 _41582_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_21141_));
 sky130_fd_sc_hd__mux2_1 _41583_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_21142_));
 sky130_fd_sc_hd__mux2_1 _41584_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_21105_));
 sky130_fd_sc_hd__mux2_1 _41585_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_21106_));
 sky130_fd_sc_hd__mux2_1 _41586_ (.A0(_00271_),
    .A1(_00216_),
    .S(net513),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _41587_ (.A0(_00265_),
    .A1(_00216_),
    .S(net513),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _41588_ (.A0(_00259_),
    .A1(_00216_),
    .S(net513),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _41589_ (.A0(_00253_),
    .A1(_00216_),
    .S(net513),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _41590_ (.A0(_00247_),
    .A1(_00216_),
    .S(net513),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _41591_ (.A0(_00233_),
    .A1(_00216_),
    .S(net513),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _41592_ (.A0(_00219_),
    .A1(_00216_),
    .S(net513),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _41593_ (.A0(_00188_),
    .A1(_00216_),
    .S(net513),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _41594_ (.A0(_00270_),
    .A1(_00271_),
    .S(net513),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _41595_ (.A0(_00246_),
    .A1(_00216_),
    .S(net514),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _41596_ (.A0(_00243_),
    .A1(_00245_),
    .S(net514),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _41597_ (.A0(_00239_),
    .A1(_00242_),
    .S(net514),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _41598_ (.A0(_00264_),
    .A1(_00265_),
    .S(net513),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _41599_ (.A0(_00232_),
    .A1(_00216_),
    .S(net514),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _41600_ (.A0(_00229_),
    .A1(_00231_),
    .S(net514),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _41601_ (.A0(_00225_),
    .A1(_00228_),
    .S(net514),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _41602_ (.A0(_00258_),
    .A1(_00259_),
    .S(net513),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _41603_ (.A0(_00218_),
    .A1(_00216_),
    .S(net514),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _41604_ (.A0(_00210_),
    .A1(_00214_),
    .S(net514),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _41605_ (.A0(_00202_),
    .A1(_00207_),
    .S(net514),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _41606_ (.A0(_00252_),
    .A1(_00253_),
    .S(net513),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _41607_ (.A0(_00187_),
    .A1(_00216_),
    .S(net514),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _41608_ (.A0(_00180_),
    .A1(_00184_),
    .S(net514),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _41609_ (.A0(_00172_),
    .A1(_00177_),
    .S(net514),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _41610_ (.A0(_00244_),
    .A1(_00247_),
    .S(net513),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _41611_ (.A0(_00245_),
    .A1(_00246_),
    .S(net514),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _41612_ (.A0(_00217_),
    .A1(_00216_),
    .S(net515),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _41613_ (.A0(_00213_),
    .A1(_00215_),
    .S(net515),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _41614_ (.A0(_00242_),
    .A1(_00243_),
    .S(net514),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _41615_ (.A0(_00209_),
    .A1(_00212_),
    .S(net515),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _41616_ (.A0(_00206_),
    .A1(_00208_),
    .S(net515),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _41617_ (.A0(_00238_),
    .A1(_00239_),
    .S(net514),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _41618_ (.A0(_00201_),
    .A1(_00205_),
    .S(net515),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _41619_ (.A0(_00198_),
    .A1(_00200_),
    .S(net515),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _41620_ (.A0(_00194_),
    .A1(_00197_),
    .S(net515),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _41621_ (.A0(_00230_),
    .A1(_00233_),
    .S(net513),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _41622_ (.A0(_00231_),
    .A1(_00232_),
    .S(net514),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _41623_ (.A0(_00186_),
    .A1(_00216_),
    .S(net515),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _41624_ (.A0(_00183_),
    .A1(_00185_),
    .S(net515),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _41625_ (.A0(_00228_),
    .A1(_00229_),
    .S(net514),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _41626_ (.A0(_00179_),
    .A1(_00182_),
    .S(net515),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _41627_ (.A0(_00176_),
    .A1(_00178_),
    .S(net515),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _41628_ (.A0(_00224_),
    .A1(_00225_),
    .S(net514),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _41629_ (.A0(_00171_),
    .A1(_00175_),
    .S(net515),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _41630_ (.A0(_00168_),
    .A1(_00170_),
    .S(net515),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _41631_ (.A0(_00164_),
    .A1(_00167_),
    .S(net515),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _41632_ (.A0(_00211_),
    .A1(_00219_),
    .S(net513),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _41633_ (.A0(_00214_),
    .A1(_00218_),
    .S(net514),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _41634_ (.A0(_00215_),
    .A1(_00217_),
    .S(net515),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _41635_ (.A0(net330),
    .A1(_00216_),
    .S(net516),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _41636_ (.A0(net327),
    .A1(net329),
    .S(net516),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _41637_ (.A0(_00212_),
    .A1(_00213_),
    .S(net515),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _41638_ (.A0(net325),
    .A1(net326),
    .S(net516),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _41639_ (.A0(net323),
    .A1(net324),
    .S(net516),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _41640_ (.A0(_00207_),
    .A1(_00210_),
    .S(net514),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _41641_ (.A0(_00208_),
    .A1(_00209_),
    .S(net515),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _41642_ (.A0(net321),
    .A1(net322),
    .S(net516),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _41643_ (.A0(net319),
    .A1(net320),
    .S(net516),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _41644_ (.A0(_00205_),
    .A1(_00206_),
    .S(net515),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _41645_ (.A0(net316),
    .A1(net318),
    .S(net516),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _41646_ (.A0(net314),
    .A1(net315),
    .S(net516),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _41647_ (.A0(_00199_),
    .A1(_00202_),
    .S(net514),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _41648_ (.A0(_00200_),
    .A1(_00201_),
    .S(net515),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _41649_ (.A0(net312),
    .A1(net313),
    .S(net516),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _41650_ (.A0(net310),
    .A1(net311),
    .S(net516),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _41651_ (.A0(_00197_),
    .A1(_00198_),
    .S(net515),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _41652_ (.A0(net308),
    .A1(net309),
    .S(net516),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _41653_ (.A0(net337),
    .A1(net307),
    .S(net516),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _41654_ (.A0(_00193_),
    .A1(_00194_),
    .S(net515),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _41655_ (.A0(net335),
    .A1(net336),
    .S(net516),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _41656_ (.A0(net333),
    .A1(net334),
    .S(net516),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _41657_ (.A0(net331),
    .A1(net332),
    .S(net516),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _41658_ (.A0(_00181_),
    .A1(_00188_),
    .S(net513),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _41659_ (.A0(_00184_),
    .A1(_00187_),
    .S(net514),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _41660_ (.A0(_00185_),
    .A1(_00186_),
    .S(net515),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _41661_ (.A0(net329),
    .A1(net330),
    .S(net516),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _41662_ (.A0(net326),
    .A1(net327),
    .S(net516),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _41663_ (.A0(_00182_),
    .A1(_00183_),
    .S(net515),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _41664_ (.A0(net324),
    .A1(net325),
    .S(net516),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _41665_ (.A0(net322),
    .A1(net323),
    .S(net516),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _41666_ (.A0(_00177_),
    .A1(_00180_),
    .S(net514),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _41667_ (.A0(_00178_),
    .A1(_00179_),
    .S(net515),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _41668_ (.A0(net320),
    .A1(net321),
    .S(net516),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _41669_ (.A0(net318),
    .A1(net319),
    .S(net516),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _41670_ (.A0(_00175_),
    .A1(_00176_),
    .S(net515),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _41671_ (.A0(net315),
    .A1(net316),
    .S(net516),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _41672_ (.A0(net313),
    .A1(net314),
    .S(net516),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _41673_ (.A0(_00169_),
    .A1(_00172_),
    .S(net514),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _41674_ (.A0(_00170_),
    .A1(_00171_),
    .S(net515),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _41675_ (.A0(net311),
    .A1(net312),
    .S(net516),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _41676_ (.A0(net309),
    .A1(net310),
    .S(net516),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _41677_ (.A0(_00167_),
    .A1(_00168_),
    .S(net515),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _41678_ (.A0(net307),
    .A1(net308),
    .S(net516),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _41679_ (.A0(net336),
    .A1(net337),
    .S(net516),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _41680_ (.A0(_00163_),
    .A1(_00164_),
    .S(net515),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _41681_ (.A0(net334),
    .A1(net335),
    .S(net516),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _41682_ (.A0(net332),
    .A1(net333),
    .S(net516),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _41683_ (.A0(net328),
    .A1(net331),
    .S(net516),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _41684_ (.A0(net327),
    .A1(net326),
    .S(net516),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _41685_ (.A0(net326),
    .A1(net325),
    .S(net200),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _41686_ (.A0(_00140_),
    .A1(_00132_),
    .S(net515),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _41687_ (.A0(net325),
    .A1(net324),
    .S(net516),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _41688_ (.A0(_00136_),
    .A1(_00128_),
    .S(net211),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _41689_ (.A0(net324),
    .A1(net323),
    .S(net516),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _41690_ (.A0(_00132_),
    .A1(_00123_),
    .S(net515),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _41691_ (.A0(net323),
    .A1(net322),
    .S(net516),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _41692_ (.A0(_00128_),
    .A1(_00117_),
    .S(net211),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _41693_ (.A0(net322),
    .A1(net321),
    .S(net516),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _41694_ (.A0(_00098_),
    .A1(_00100_),
    .S(net514),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _41695_ (.A0(_00124_),
    .A1(_00097_),
    .S(net514),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _41696_ (.A0(_00123_),
    .A1(_00111_),
    .S(net515),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _41697_ (.A0(net321),
    .A1(net320),
    .S(net516),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _41698_ (.A0(_00101_),
    .A1(_00094_),
    .S(net222),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _41699_ (.A0(_00088_),
    .A1(_00090_),
    .S(net222),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _41700_ (.A0(_00118_),
    .A1(_00087_),
    .S(net222),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _41701_ (.A0(_00117_),
    .A1(_00105_),
    .S(net211),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _41702_ (.A0(net320),
    .A1(net319),
    .S(net200),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _41703_ (.A0(_00091_),
    .A1(_00084_),
    .S(net222),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _41704_ (.A0(_00074_),
    .A1(_00078_),
    .S(net514),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _41705_ (.A0(_00112_),
    .A1(_00071_),
    .S(net514),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _41706_ (.A0(_00111_),
    .A1(_00096_),
    .S(net515),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _41707_ (.A0(net319),
    .A1(net318),
    .S(net516),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _41708_ (.A0(_00081_),
    .A1(_00067_),
    .S(net222),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _41709_ (.A0(_00056_),
    .A1(_00060_),
    .S(net222),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _41710_ (.A0(_00106_),
    .A1(_00053_),
    .S(net222),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _41711_ (.A0(_00105_),
    .A1(_00086_),
    .S(net211),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _41712_ (.A0(net318),
    .A1(net316),
    .S(net200),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _41713_ (.A0(_00063_),
    .A1(_00049_),
    .S(net222),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _41714_ (.A0(_00100_),
    .A1(_00101_),
    .S(net514),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _41715_ (.A0(_00077_),
    .A1(_00079_),
    .S(net515),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _41716_ (.A0(_00073_),
    .A1(_00076_),
    .S(net515),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _41717_ (.A0(_00097_),
    .A1(_00098_),
    .S(net514),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _41718_ (.A0(_00070_),
    .A1(_00072_),
    .S(net515),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _41719_ (.A0(_00096_),
    .A1(_00069_),
    .S(net515),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _41720_ (.A0(net316),
    .A1(net315),
    .S(net516),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_2 _41721_ (.A0(_00080_),
    .A1(_00066_),
    .S(net515),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _41722_ (.A0(_00090_),
    .A1(_00091_),
    .S(net222),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _41723_ (.A0(_00059_),
    .A1(_00061_),
    .S(net211),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _41724_ (.A0(_00055_),
    .A1(_00058_),
    .S(net211),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _41725_ (.A0(_00087_),
    .A1(_00088_),
    .S(net222),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _41726_ (.A0(_00052_),
    .A1(_00054_),
    .S(net211),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _41727_ (.A0(_00086_),
    .A1(_00051_),
    .S(net211),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _41728_ (.A0(net315),
    .A1(net314),
    .S(net200),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_2 _41729_ (.A0(_00062_),
    .A1(_00048_),
    .S(net211),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _41730_ (.A0(_00078_),
    .A1(_00081_),
    .S(net222),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _41731_ (.A0(_00079_),
    .A1(_00080_),
    .S(net515),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _41732_ (.A0(net331),
    .A1(net328),
    .S(net200),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _41733_ (.A0(net333),
    .A1(net332),
    .S(net200),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _41734_ (.A0(_00076_),
    .A1(_00077_),
    .S(net515),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _41735_ (.A0(net335),
    .A1(net334),
    .S(net200),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _41736_ (.A0(net337),
    .A1(net336),
    .S(net200),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _41737_ (.A0(_00071_),
    .A1(_00074_),
    .S(net514),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _41738_ (.A0(_00072_),
    .A1(_00073_),
    .S(net515),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _41739_ (.A0(net308),
    .A1(net307),
    .S(net200),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _41740_ (.A0(net310),
    .A1(net309),
    .S(net200),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _41741_ (.A0(_00069_),
    .A1(_00070_),
    .S(net515),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _41742_ (.A0(net312),
    .A1(net311),
    .S(net516),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _41743_ (.A0(net314),
    .A1(net313),
    .S(net516),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _41744_ (.A0(net317),
    .A1(net306),
    .S(net200),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _41745_ (.A0(_00060_),
    .A1(_00063_),
    .S(net222),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _41746_ (.A0(_00061_),
    .A1(_00062_),
    .S(net211),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _41747_ (.A0(net328),
    .A1(net317),
    .S(net200),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _41748_ (.A0(net332),
    .A1(net331),
    .S(net200),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _41749_ (.A0(_00058_),
    .A1(_00059_),
    .S(net211),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _41750_ (.A0(net334),
    .A1(net333),
    .S(net200),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _41751_ (.A0(net336),
    .A1(net335),
    .S(net200),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _41752_ (.A0(_00053_),
    .A1(_00056_),
    .S(net222),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _41753_ (.A0(_00054_),
    .A1(_00055_),
    .S(net211),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _41754_ (.A0(net307),
    .A1(net337),
    .S(net200),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _41755_ (.A0(net309),
    .A1(net308),
    .S(net200),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _41756_ (.A0(_00051_),
    .A1(_00052_),
    .S(net211),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _41757_ (.A0(net311),
    .A1(net310),
    .S(net200),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _41758_ (.A0(net313),
    .A1(net312),
    .S(net200),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _41759_ (.A0(_02408_),
    .A1(net362),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _41760_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_2 _41761_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _41762_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _41763_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _41764_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _41765_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _41766_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _41767_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _41768_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _41769_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _41770_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _41771_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _41772_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _41773_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _41774_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _41775_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _41776_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _41777_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _41778_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _41779_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _41780_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _41781_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _41782_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _41783_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _41784_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _41785_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _41786_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _41787_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _41788_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _41789_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _41790_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _41791_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _41792_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _41793_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _41794_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _41795_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(_01208_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _41796_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _41797_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _41798_ (.A0(_02056_),
    .A1(_02055_),
    .S(_01714_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_2 _41799_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _41800_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _41801_ (.A0(_01908_),
    .A1(_02052_),
    .S(_01816_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _41802_ (.A0(_02047_),
    .A1(_02046_),
    .S(_01714_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_2 _41803_ (.A0(_02049_),
    .A1(_02048_),
    .S(_01717_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _41804_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _41805_ (.A0(_01908_),
    .A1(_02043_),
    .S(_01816_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_2 _41806_ (.A0(_02038_),
    .A1(_02037_),
    .S(_01714_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _41807_ (.A0(_02040_),
    .A1(_02039_),
    .S(_01717_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _41808_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _41809_ (.A0(_01908_),
    .A1(_02034_),
    .S(_01816_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_2 _41810_ (.A0(_02029_),
    .A1(_02028_),
    .S(_01714_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_2 _41811_ (.A0(_02031_),
    .A1(_02030_),
    .S(_01717_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _41812_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_2 _41813_ (.A0(_01908_),
    .A1(_02025_),
    .S(_01816_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_2 _41814_ (.A0(_02020_),
    .A1(_02019_),
    .S(_01714_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_2 _41815_ (.A0(_02022_),
    .A1(_02021_),
    .S(_01717_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _41816_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _41817_ (.A0(_01908_),
    .A1(_02016_),
    .S(_01816_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_2 _41818_ (.A0(_02011_),
    .A1(_02010_),
    .S(_01714_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _41819_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _41820_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_2 _41821_ (.A0(_01908_),
    .A1(_02007_),
    .S(_01816_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_2 _41822_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_2 _41823_ (.A0(_02004_),
    .A1(_02003_),
    .S(_01717_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _41824_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_2 _41825_ (.A0(_01908_),
    .A1(_01998_),
    .S(net506),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _41826_ (.A0(_01993_),
    .A1(_01992_),
    .S(_01714_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_2 _41827_ (.A0(_01995_),
    .A1(_01994_),
    .S(_01717_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _41828_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(net519),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _41829_ (.A0(_01908_),
    .A1(_01989_),
    .S(_01816_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_2 _41830_ (.A0(_01984_),
    .A1(_01983_),
    .S(_01714_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_2 _41831_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _41832_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(net519),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _41833_ (.A0(_01908_),
    .A1(_01980_),
    .S(_01816_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _41834_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _41835_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _41836_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(net519),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _41837_ (.A0(_01908_),
    .A1(_01971_),
    .S(net506),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_2 _41838_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_2 _41839_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _41840_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(net519),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _41841_ (.A0(_01908_),
    .A1(_01962_),
    .S(net506),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _41842_ (.A0(_01957_),
    .A1(_01956_),
    .S(_01714_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_2 _41843_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _41844_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(net519),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _41845_ (.A0(_01908_),
    .A1(_01953_),
    .S(net506),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _41846_ (.A0(_01948_),
    .A1(_01947_),
    .S(_01714_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_2 _41847_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _41848_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _41849_ (.A0(_01908_),
    .A1(_01944_),
    .S(net506),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _41850_ (.A0(_01939_),
    .A1(_01938_),
    .S(_01714_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_2 _41851_ (.A0(_01941_),
    .A1(_01940_),
    .S(_01717_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _41852_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(net519),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _41853_ (.A0(_01908_),
    .A1(_01935_),
    .S(net506),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_2 _41854_ (.A0(_01930_),
    .A1(_01929_),
    .S(_01714_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_2 _41855_ (.A0(_01932_),
    .A1(_01931_),
    .S(_01717_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _41856_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(net519),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _41857_ (.A0(_01908_),
    .A1(_01926_),
    .S(net506),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_2 _41858_ (.A0(_01921_),
    .A1(_01920_),
    .S(_01714_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_2 _41859_ (.A0(_01923_),
    .A1(_01922_),
    .S(_01717_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_2 _41860_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(net519),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _41861_ (.A0(_01908_),
    .A1(_01917_),
    .S(net506),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_2 _41862_ (.A0(_01912_),
    .A1(_01911_),
    .S(_01714_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_2 _41863_ (.A0(_01914_),
    .A1(_01913_),
    .S(_01717_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_2 _41864_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(net519),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_2 _41865_ (.A0(_01908_),
    .A1(_01907_),
    .S(net506),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _41866_ (.A0(_01906_),
    .A1(_01904_),
    .S(net450),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _41867_ (.A0(net527),
    .A1(net57),
    .S(net317),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _41868_ (.A0(_01899_),
    .A1(_01898_),
    .S(_01714_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_2 _41869_ (.A0(_01901_),
    .A1(_01900_),
    .S(_01717_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_2 _41870_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(net519),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _41871_ (.A0(_01895_),
    .A1(_01894_),
    .S(net506),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _41872_ (.A0(_01893_),
    .A1(_01891_),
    .S(net450),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _41873_ (.A0(net38),
    .A1(net523),
    .S(net317),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _41874_ (.A0(_01886_),
    .A1(_01885_),
    .S(_01714_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_2 _41875_ (.A0(_01888_),
    .A1(_01887_),
    .S(_01717_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_4 _41876_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(net519),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _41877_ (.A0(_01882_),
    .A1(_01881_),
    .S(net506),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _41878_ (.A0(_01880_),
    .A1(_01878_),
    .S(net451),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _41879_ (.A0(net37),
    .A1(net54),
    .S(net317),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _41880_ (.A0(_01873_),
    .A1(_01872_),
    .S(_01714_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_2 _41881_ (.A0(_01875_),
    .A1(_01874_),
    .S(_01717_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_4 _41882_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(net519),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_2 _41883_ (.A0(_01869_),
    .A1(_01868_),
    .S(net506),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _41884_ (.A0(_01867_),
    .A1(_01865_),
    .S(net450),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _41885_ (.A0(net528),
    .A1(net53),
    .S(net317),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_2 _41886_ (.A0(_01860_),
    .A1(_01859_),
    .S(_01714_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_2 _41887_ (.A0(_01862_),
    .A1(_01861_),
    .S(_01717_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_4 _41888_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(net519),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _41889_ (.A0(_01856_),
    .A1(_01855_),
    .S(net506),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _41890_ (.A0(_01854_),
    .A1(_01852_),
    .S(net451),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _41891_ (.A0(net35),
    .A1(net52),
    .S(net317),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _41892_ (.A0(_01847_),
    .A1(_01846_),
    .S(_01714_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_2 _41893_ (.A0(_01849_),
    .A1(_01848_),
    .S(_01717_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_4 _41894_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(net519),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_2 _41895_ (.A0(_01843_),
    .A1(_01842_),
    .S(net506),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _41896_ (.A0(_01841_),
    .A1(_01839_),
    .S(net450),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _41897_ (.A0(net34),
    .A1(net51),
    .S(net317),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_2 _41898_ (.A0(_01834_),
    .A1(_01833_),
    .S(_01714_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_2 _41899_ (.A0(_01836_),
    .A1(_01835_),
    .S(_01717_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_4 _41900_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(net519),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _41901_ (.A0(_01830_),
    .A1(_01829_),
    .S(net506),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _41902_ (.A0(_01828_),
    .A1(_01826_),
    .S(net451),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _41903_ (.A0(net64),
    .A1(net50),
    .S(net317),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _41904_ (.A0(_01821_),
    .A1(_01820_),
    .S(_01714_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_2 _41905_ (.A0(_01823_),
    .A1(_01822_),
    .S(_01717_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_4 _41906_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(net519),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _41907_ (.A0(_01817_),
    .A1(_01815_),
    .S(net506),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _41908_ (.A0(_01814_),
    .A1(_01812_),
    .S(net450),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _41909_ (.A0(net63),
    .A1(net49),
    .S(net317),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_2 _41910_ (.A0(_01807_),
    .A1(_01806_),
    .S(_01714_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_2 _41911_ (.A0(_01809_),
    .A1(_01808_),
    .S(_01717_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_8 _41912_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(net519),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _41913_ (.A0(_01803_),
    .A1(_01799_),
    .S(net450),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _41914_ (.A0(net62),
    .A1(net48),
    .S(net317),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _41915_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _41916_ (.A0(_01794_),
    .A1(_01793_),
    .S(_01714_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_2 _41917_ (.A0(_01796_),
    .A1(_01795_),
    .S(_01717_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_8 _41918_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(net519),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_2 _41919_ (.A0(_01790_),
    .A1(_01786_),
    .S(net450),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _41920_ (.A0(net61),
    .A1(net47),
    .S(net317),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _41921_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _41922_ (.A0(_01781_),
    .A1(_01780_),
    .S(_01714_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_2 _41923_ (.A0(_01783_),
    .A1(_01782_),
    .S(_01717_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_8 _41924_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(net519),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _41925_ (.A0(_01777_),
    .A1(_01773_),
    .S(net451),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _41926_ (.A0(net522),
    .A1(net46),
    .S(net317),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _41927_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _41928_ (.A0(_01768_),
    .A1(_01767_),
    .S(_01714_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_2 _41929_ (.A0(_01770_),
    .A1(_01769_),
    .S(_01717_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_8 _41930_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(net519),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _41931_ (.A0(_01764_),
    .A1(_01760_),
    .S(net450),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _41932_ (.A0(net59),
    .A1(net524),
    .S(net317),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _41933_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _41934_ (.A0(_01755_),
    .A1(_01754_),
    .S(_01714_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_2 _41935_ (.A0(_01757_),
    .A1(_01756_),
    .S(_01717_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_4 _41936_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(net519),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _41937_ (.A0(_01751_),
    .A1(_01747_),
    .S(net450),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _41938_ (.A0(net58),
    .A1(net526),
    .S(net317),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _41939_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _41940_ (.A0(_01742_),
    .A1(_01741_),
    .S(_01714_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_2 _41941_ (.A0(_01744_),
    .A1(_01743_),
    .S(_01717_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_4 _41942_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(net519),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _41943_ (.A0(_01738_),
    .A1(_01734_),
    .S(net450),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _41944_ (.A0(net55),
    .A1(net42),
    .S(net317),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _41945_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _41946_ (.A0(_01729_),
    .A1(_01728_),
    .S(_01714_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_2 _41947_ (.A0(_01731_),
    .A1(_01730_),
    .S(_01717_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_2 _41948_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(net519),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _41949_ (.A0(_01725_),
    .A1(_01721_),
    .S(net450),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _41950_ (.A0(net525),
    .A1(net41),
    .S(net317),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _41951_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _41952_ (.A0(_01715_),
    .A1(_02559_),
    .S(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _41953_ (.A0(_01718_),
    .A1(_01716_),
    .S(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_2 _41954_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(net519),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _41955_ (.A0(_01711_),
    .A1(_01707_),
    .S(net450),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _41956_ (.A0(net33),
    .A1(net40),
    .S(net317),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _41957_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _41958_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _41959_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _41960_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _41961_ (.A0(_01693_),
    .A1(net273),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _41962_ (.A0(_01690_),
    .A1(net272),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _41963_ (.A0(_01687_),
    .A1(net271),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _41964_ (.A0(_01684_),
    .A1(net270),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _41965_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(net511),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _41966_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _41967_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(net511),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _41968_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _41969_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(net511),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _41970_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _41971_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(net511),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _41972_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _41973_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(net511),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _41974_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _41975_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(net511),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _41976_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _41977_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(net511),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _41978_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _41979_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(net511),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _41980_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _41981_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(net511),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _41982_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _41983_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(net511),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _41984_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _41985_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(net511),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _41986_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _41987_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(net511),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _41988_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _41989_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(net511),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _41990_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _41991_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(net511),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _41992_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _41993_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(net511),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _41994_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _41995_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(net511),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_2 _41996_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _41997_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(net511),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _41998_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _41999_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(net511),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _42000_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _42001_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(net511),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _42002_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _42003_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(net511),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _42004_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _42005_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(net511),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _42006_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _42007_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(net511),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _42008_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _42009_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(net511),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _42010_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _42011_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(net511),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _42012_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _42013_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(net511),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _42014_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _42015_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(net511),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _42016_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _42017_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(net511),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _42018_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_2 _42019_ (.A0(_01474_),
    .A1(_01471_),
    .S(net472),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _42020_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(net511),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _42021_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _42022_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(net511),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _42023_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _42024_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(net511),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _42025_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _42026_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _42027_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _42028_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(net410),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _42029_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(net410),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _42030_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(net410),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _42031_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(net410),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _42032_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(net410),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _42033_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(net410),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _42034_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(net410),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _42035_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(net410),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _42036_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(net410),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _42037_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(net410),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _42038_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(net410),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _42039_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(net410),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _42040_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(net410),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _42041_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(net410),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _42042_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(net410),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _42043_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(_01208_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _42044_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(_01208_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _42045_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(_01208_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _42046_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(net410),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _42047_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(net410),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _42048_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(_01208_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _42049_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(_01208_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _42050_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(_01208_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _42051_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(_01208_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _42052_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(_01208_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _42053_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(_01208_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _42054_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(_01208_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _42055_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(_01208_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _42056_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(_01208_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_2 _42057_ (.A0(_01206_),
    .A1(_01201_),
    .S(net462),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_4 _42058_ (.A0(_01179_),
    .A1(_01174_),
    .S(_00368_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_4 _42059_ (.A0(_01152_),
    .A1(_01147_),
    .S(_00368_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_4 _42060_ (.A0(_01125_),
    .A1(_01120_),
    .S(_00368_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_4 _42061_ (.A0(_01098_),
    .A1(_01093_),
    .S(_00368_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_2 _42062_ (.A0(_01071_),
    .A1(_01066_),
    .S(net462),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_4 _42063_ (.A0(_01044_),
    .A1(_01039_),
    .S(net461),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_4 _42064_ (.A0(_01017_),
    .A1(_01012_),
    .S(net461),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_4 _42065_ (.A0(_00990_),
    .A1(_00985_),
    .S(net461),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_8 _42066_ (.A0(_00963_),
    .A1(_00958_),
    .S(net461),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_8 _42067_ (.A0(_00936_),
    .A1(_00931_),
    .S(net462),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_4 _42068_ (.A0(_00909_),
    .A1(_00904_),
    .S(net461),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_4 _42069_ (.A0(_00882_),
    .A1(_00877_),
    .S(net462),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_4 _42070_ (.A0(_00855_),
    .A1(_00850_),
    .S(net462),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_4 _42071_ (.A0(_00828_),
    .A1(_00823_),
    .S(net462),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_4 _42072_ (.A0(_00801_),
    .A1(_00796_),
    .S(net462),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_4 _42073_ (.A0(_00774_),
    .A1(_00769_),
    .S(net462),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_4 _42074_ (.A0(_00747_),
    .A1(_00742_),
    .S(net462),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_4 _42075_ (.A0(_00720_),
    .A1(_00715_),
    .S(net460),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_8 _42076_ (.A0(_00693_),
    .A1(_00688_),
    .S(net460),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_8 _42077_ (.A0(_00666_),
    .A1(_00661_),
    .S(net460),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_8 _42078_ (.A0(_00639_),
    .A1(_00634_),
    .S(net460),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_8 _42079_ (.A0(_00612_),
    .A1(_00607_),
    .S(net460),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_4 _42080_ (.A0(_00585_),
    .A1(_00580_),
    .S(net460),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_8 _42081_ (.A0(_00558_),
    .A1(_00553_),
    .S(net460),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_8 _42082_ (.A0(_00531_),
    .A1(_00526_),
    .S(net461),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_8 _42083_ (.A0(_00504_),
    .A1(_00499_),
    .S(net460),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_8 _42084_ (.A0(_00477_),
    .A1(_00472_),
    .S(net460),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_8 _42085_ (.A0(_00450_),
    .A1(_00445_),
    .S(net461),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_8 _42086_ (.A0(_00423_),
    .A1(_00418_),
    .S(net461),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_4 _42087_ (.A0(_00396_),
    .A1(_00391_),
    .S(net461),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_2 _42088_ (.A0(_00369_),
    .A1(_00365_),
    .S(net462),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_8 _42089_ (.A0(_00366_),
    .A1(_00367_),
    .S(\cpu_state[3] ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_8 _42090_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(net517),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_4 _42091_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(net517),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_4 _42092_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(\cpu_state[3] ),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_8 _42093_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(net517),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _42094_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _42095_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _42096_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _42097_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _42098_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _42099_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_4 _42100_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _42101_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _42102_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _42103_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _42104_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _42105_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_2 _42106_ (.A0(\mem_rdata_q[6] ),
    .A1(net61),
    .S(net437),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_4 _42107_ (.A0(\mem_rdata_q[5] ),
    .A1(net522),
    .S(net437),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_4 _42108_ (.A0(\mem_rdata_q[4] ),
    .A1(net59),
    .S(net437),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_2 _42109_ (.A0(\mem_rdata_q[3] ),
    .A1(net58),
    .S(net437),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _42110_ (.A0(\mem_rdata_q[2] ),
    .A1(net55),
    .S(net437),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _42111_ (.A0(\mem_rdata_q[1] ),
    .A1(net525),
    .S(net437),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _42112_ (.A0(\mem_rdata_q[0] ),
    .A1(net33),
    .S(net437),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _42113_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(net518),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _42114_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _42115_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _42116_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _42117_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _42118_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(net511),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _42119_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _42120_ (.A0(_00126_),
    .A1(_00122_),
    .S(net513),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _42121_ (.A0(_00120_),
    .A1(_00116_),
    .S(net225),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _42122_ (.A0(_00114_),
    .A1(_00110_),
    .S(net513),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _42123_ (.A0(_00108_),
    .A1(_00104_),
    .S(net225),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _42124_ (.A0(_00102_),
    .A1(_00095_),
    .S(net513),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _42125_ (.A0(_00092_),
    .A1(_00085_),
    .S(net225),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_2 _42126_ (.A0(_00082_),
    .A1(_00068_),
    .S(net513),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _42127_ (.A0(_00064_),
    .A1(_00050_),
    .S(net225),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _42128_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _42129_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _42130_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _42131_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _42132_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_2 _42133_ (.A0(_01682_),
    .A1(_02581_),
    .S(net415),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _42134_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _42135_ (.A0(_01678_),
    .A1(_02580_),
    .S(net415),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _42136_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _42137_ (.A0(_01674_),
    .A1(_02579_),
    .S(net415),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _42138_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _42139_ (.A0(_01670_),
    .A1(_02578_),
    .S(net415),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _42140_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _42141_ (.A0(_01666_),
    .A1(_02577_),
    .S(net414),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _42142_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _42143_ (.A0(_01662_),
    .A1(_02576_),
    .S(net414),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _42144_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _42145_ (.A0(_01658_),
    .A1(_02575_),
    .S(net414),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _42146_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _42147_ (.A0(_01654_),
    .A1(_02574_),
    .S(net414),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _42148_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _42149_ (.A0(_01650_),
    .A1(_02573_),
    .S(net414),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _42150_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _42151_ (.A0(_01646_),
    .A1(_02572_),
    .S(net414),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _42152_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _42153_ (.A0(_01642_),
    .A1(_02570_),
    .S(net414),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _42154_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _42155_ (.A0(_01638_),
    .A1(_02569_),
    .S(net414),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _42156_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _42157_ (.A0(_01634_),
    .A1(_02568_),
    .S(net414),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _42158_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _42159_ (.A0(_01630_),
    .A1(_02567_),
    .S(net414),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _42160_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _42161_ (.A0(_01626_),
    .A1(_02566_),
    .S(net414),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _42162_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _42163_ (.A0(_01622_),
    .A1(_02565_),
    .S(net414),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _42164_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _42165_ (.A0(_01618_),
    .A1(_02564_),
    .S(net414),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _42166_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _42167_ (.A0(_01614_),
    .A1(_02563_),
    .S(net415),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _42168_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _42169_ (.A0(_01610_),
    .A1(_02562_),
    .S(net415),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _42170_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _42171_ (.A0(_01606_),
    .A1(_02561_),
    .S(net415),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _42172_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _42173_ (.A0(_01602_),
    .A1(_02589_),
    .S(net415),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _42174_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _42175_ (.A0(_01598_),
    .A1(_02588_),
    .S(net415),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _42176_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _42177_ (.A0(_01594_),
    .A1(_02587_),
    .S(net415),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _42178_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _42179_ (.A0(_01590_),
    .A1(_02586_),
    .S(net415),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _42180_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _42181_ (.A0(_01586_),
    .A1(_02585_),
    .S(net415),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _42182_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _42183_ (.A0(_01582_),
    .A1(_02584_),
    .S(_00308_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _42184_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _42185_ (.A0(_01578_),
    .A1(_02583_),
    .S(net415),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _42186_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _42187_ (.A0(_01574_),
    .A1(_02582_),
    .S(_00308_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _42188_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _42189_ (.A0(_01570_),
    .A1(_02571_),
    .S(_00308_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _42190_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _42191_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _42192_ (.A0(_01564_),
    .A1(_01565_),
    .S(net459),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _42193_ (.A0(_01566_),
    .A1(_02560_),
    .S(_00308_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _42194_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _42195_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _42196_ (.A0(_01559_),
    .A1(_02590_),
    .S(net459),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _42197_ (.A0(_01560_),
    .A1(_02590_),
    .S(_00308_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _42198_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _42199_ (.A0(_01464_),
    .A1(_01463_),
    .S(net509),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _42200_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _42201_ (.A0(_01461_),
    .A1(_01460_),
    .S(net509),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _42202_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _42203_ (.A0(_01458_),
    .A1(_01457_),
    .S(net509),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _42204_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _42205_ (.A0(_01455_),
    .A1(_01454_),
    .S(net509),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _42206_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _42207_ (.A0(_01452_),
    .A1(_01451_),
    .S(net509),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _42208_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _42209_ (.A0(_01449_),
    .A1(_01448_),
    .S(net509),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _42210_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _42211_ (.A0(_01446_),
    .A1(_01445_),
    .S(net509),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _42212_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _42213_ (.A0(_01443_),
    .A1(_01442_),
    .S(net509),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _42214_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _42215_ (.A0(_01440_),
    .A1(_01439_),
    .S(net509),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _42216_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _42217_ (.A0(_01437_),
    .A1(_01436_),
    .S(net509),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _42218_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _42219_ (.A0(_01434_),
    .A1(_01433_),
    .S(net509),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _42220_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _42221_ (.A0(_01431_),
    .A1(_01430_),
    .S(net509),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _42222_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _42223_ (.A0(_01428_),
    .A1(_01427_),
    .S(net509),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _42224_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _42225_ (.A0(_01425_),
    .A1(_01424_),
    .S(net509),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _42226_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _42227_ (.A0(_01422_),
    .A1(_01421_),
    .S(net509),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _42228_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _42229_ (.A0(_01419_),
    .A1(_01418_),
    .S(net509),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _42230_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _42231_ (.A0(_01416_),
    .A1(_01415_),
    .S(net509),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _42232_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _42233_ (.A0(_01413_),
    .A1(_01412_),
    .S(net510),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _42234_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _42235_ (.A0(_01410_),
    .A1(_01409_),
    .S(net510),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _42236_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _42237_ (.A0(_01407_),
    .A1(_01406_),
    .S(net510),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _42238_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _42239_ (.A0(_01404_),
    .A1(_01403_),
    .S(net510),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _42240_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _42241_ (.A0(_01401_),
    .A1(_01400_),
    .S(net510),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _42242_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _42243_ (.A0(_01398_),
    .A1(_01397_),
    .S(net510),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _42244_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _42245_ (.A0(_01395_),
    .A1(_01394_),
    .S(net510),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _42246_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _42247_ (.A0(_01392_),
    .A1(_01391_),
    .S(net510),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _42248_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _42249_ (.A0(_01389_),
    .A1(_01388_),
    .S(net510),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _42250_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _42251_ (.A0(_01386_),
    .A1(_01385_),
    .S(net510),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _42252_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _42253_ (.A0(_01383_),
    .A1(_01382_),
    .S(net510),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _42254_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _42255_ (.A0(_01380_),
    .A1(_01379_),
    .S(net510),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _42256_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _42257_ (.A0(_01377_),
    .A1(_01376_),
    .S(net510),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _42258_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _42259_ (.A0(_01374_),
    .A1(_01373_),
    .S(net510),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _42260_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _42261_ (.A0(_01371_),
    .A1(_01370_),
    .S(net510),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _42262_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(net508),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _42263_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(net517),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _42264_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(net507),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _42265_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(net517),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _42266_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(net507),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_2 _42267_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(net517),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _42268_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(net507),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _42269_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(net517),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _42270_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(net507),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _42271_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(net517),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _42272_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(net507),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _42273_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(net517),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _42274_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(net507),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _42275_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(net517),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _42276_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(net507),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _42277_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(net517),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _42278_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(net507),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _42279_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(net517),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _42280_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(net507),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _42281_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(net517),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _42282_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(net507),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _42283_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(net517),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _42284_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(net507),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _42285_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(net517),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _42286_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(net507),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _42287_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(net517),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _42288_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(net507),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _42289_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(net517),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _42290_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(net507),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _42291_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(net517),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _42292_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(net507),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _42293_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(net517),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _42294_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(net507),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _42295_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(net517),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _42296_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(net507),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _42297_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(net517),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _42298_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(net508),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _42299_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(net517),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _42300_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(net508),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _42301_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(net517),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _42302_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(net508),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _42303_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(net517),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _42304_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(net508),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _42305_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(net517),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _42306_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(net508),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _42307_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(net517),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _42308_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(net508),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _42309_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(net517),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _42310_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(net508),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _42311_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(net517),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _42312_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(net508),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _42313_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(net517),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _42314_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(net508),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _42315_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(net517),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _42316_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _42317_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(net508),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _42318_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(net517),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _42319_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _42320_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(net508),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _42321_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(net517),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _42322_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _42323_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(net508),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _42324_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(net517),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _42325_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _42326_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(net508),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _42327_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(net517),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _42328_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _42329_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(net508),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _42330_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(net517),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _42331_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(instr_timer),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _42332_ (.A0(_01302_),
    .A1(_01303_),
    .S(net518),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _42333_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(instr_timer),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _42334_ (.A0(_01299_),
    .A1(_01300_),
    .S(net518),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _42335_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(instr_timer),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _42336_ (.A0(_01296_),
    .A1(_01297_),
    .S(net518),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _42337_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(instr_timer),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _42338_ (.A0(_01293_),
    .A1(_01294_),
    .S(net518),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _42339_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(instr_timer),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _42340_ (.A0(_01290_),
    .A1(_01291_),
    .S(net518),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _42341_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(instr_timer),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _42342_ (.A0(_01287_),
    .A1(_01288_),
    .S(net518),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _42343_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(instr_timer),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _42344_ (.A0(_01284_),
    .A1(_01285_),
    .S(net518),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _42345_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(instr_timer),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _42346_ (.A0(_01281_),
    .A1(_01282_),
    .S(net518),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _42347_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(instr_timer),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _42348_ (.A0(_01278_),
    .A1(_01279_),
    .S(net518),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _42349_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(instr_timer),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _42350_ (.A0(_01275_),
    .A1(_01276_),
    .S(net518),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _42351_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(instr_timer),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _42352_ (.A0(_01272_),
    .A1(_01273_),
    .S(net518),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _42353_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(instr_timer),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _42354_ (.A0(_01269_),
    .A1(_01270_),
    .S(net518),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _42355_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(instr_timer),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _42356_ (.A0(_01266_),
    .A1(_01267_),
    .S(net518),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _42357_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(instr_timer),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _42358_ (.A0(_01263_),
    .A1(_01264_),
    .S(net518),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _42359_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(instr_timer),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _42360_ (.A0(_01260_),
    .A1(_01261_),
    .S(net518),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _42361_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(instr_timer),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _42362_ (.A0(_01257_),
    .A1(_01258_),
    .S(net518),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _42363_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(instr_timer),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _42364_ (.A0(_01254_),
    .A1(_01255_),
    .S(net518),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _42365_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(instr_timer),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _42366_ (.A0(_01251_),
    .A1(_01252_),
    .S(net518),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _42367_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(instr_timer),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _42368_ (.A0(_01248_),
    .A1(_01249_),
    .S(net518),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _42369_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(instr_timer),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _42370_ (.A0(_01245_),
    .A1(_01246_),
    .S(net518),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _42371_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(instr_timer),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _42372_ (.A0(_01242_),
    .A1(_01243_),
    .S(net518),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _42373_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(instr_timer),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _42374_ (.A0(_01239_),
    .A1(_01240_),
    .S(net518),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _42375_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(instr_timer),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _42376_ (.A0(_01236_),
    .A1(_01237_),
    .S(net518),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _42377_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(instr_timer),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _42378_ (.A0(_01233_),
    .A1(_01234_),
    .S(net518),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _42379_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(instr_timer),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _42380_ (.A0(_01230_),
    .A1(_01231_),
    .S(net518),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _42381_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(instr_timer),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _42382_ (.A0(_01227_),
    .A1(_01228_),
    .S(net518),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _42383_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(instr_timer),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _42384_ (.A0(_01224_),
    .A1(_01225_),
    .S(net518),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _42385_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(instr_timer),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _42386_ (.A0(_01221_),
    .A1(_01222_),
    .S(net518),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _42387_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(instr_timer),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _42388_ (.A0(_01218_),
    .A1(_01219_),
    .S(net518),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _42389_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(instr_timer),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _42390_ (.A0(_01215_),
    .A1(_01216_),
    .S(net518),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _42391_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(instr_timer),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _42392_ (.A0(_01212_),
    .A1(_01213_),
    .S(net518),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _42393_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(instr_timer),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _42394_ (.A0(_01209_),
    .A1(_01210_),
    .S(net518),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_1 _42395_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(net478),
    .S1(net491),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_1 _42396_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(net478),
    .S1(net491),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_2 _42397_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(net478),
    .S1(net491),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_2 _42398_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(net478),
    .S1(net491),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _42399_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(net478),
    .S1(net491),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_1 _42400_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(net498),
    .S1(net502),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_1 _42401_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(net479),
    .S1(net490),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_2 _42402_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(net479),
    .S1(net490),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_2 _42403_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(net479),
    .S1(net490),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_1 _42404_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(net479),
    .S1(net490),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_2 _42405_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(net479),
    .S1(net490),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_2 _42406_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(net498),
    .S1(net502),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _42407_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(net480),
    .S1(net490),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_2 _42408_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(net480),
    .S1(net490),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_2 _42409_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(net480),
    .S1(net490),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_1 _42410_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(net480),
    .S1(net490),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_1 _42411_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(net480),
    .S1(net490),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_2 _42412_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(net498),
    .S1(net502),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_2 _42413_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(net479),
    .S1(net490),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_1 _42414_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(net479),
    .S1(net490),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_2 _42415_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(net479),
    .S1(net490),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_1 _42416_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(net479),
    .S1(net490),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_2 _42417_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(net479),
    .S1(net490),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_1 _42418_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(net498),
    .S1(net502),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _42419_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(net479),
    .S1(net490),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_2 _42420_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(net479),
    .S1(net490),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_2 _42421_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(net479),
    .S1(net490),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_2 _42422_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(net479),
    .S1(net490),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_2 _42423_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(net479),
    .S1(net490),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_2 _42424_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(net498),
    .S1(net502),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_1 _42425_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(net478),
    .S1(net491),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_1 _42426_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(net480),
    .S1(net490),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_2 _42427_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(net480),
    .S1(net490),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _42428_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(net480),
    .S1(net491),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_1 _42429_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(net480),
    .S1(net490),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_2 _42430_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(net498),
    .S1(net502),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_1 _42431_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(net487),
    .S1(net496),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_2 _42432_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(net487),
    .S1(net496),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_2 _42433_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(net487),
    .S1(net496),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_1 _42434_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(net489),
    .S1(net496),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _42435_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(net487),
    .S1(net496),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_2 _42436_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(net500),
    .S1(net501),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_1 _42437_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(net486),
    .S1(net496),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_2 _42438_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(net487),
    .S1(net495),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_2 _42439_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(net487),
    .S1(net496),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_1 _42440_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(net487),
    .S1(net496),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_2 _42441_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(net487),
    .S1(net496),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_2 _42442_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(net500),
    .S1(net501),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_1 _42443_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(net487),
    .S1(net495),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_2 _42444_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(net487),
    .S1(net495),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_2 _42445_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(net487),
    .S1(net496),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_1 _42446_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(net487),
    .S1(net496),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_2 _42447_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(net487),
    .S1(net496),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_2 _42448_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(net500),
    .S1(net501),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_2 _42449_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(_00357_),
    .S1(net497),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_2 _42450_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(net489),
    .S1(net497),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_2 _42451_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(net489),
    .S1(net497),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _42452_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(_00357_),
    .S1(net497),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_2 _42453_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(_00357_),
    .S1(net497),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_2 _42454_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(net500),
    .S1(_00362_),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_2 _42455_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(net488),
    .S1(net497),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_2 _42456_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(net488),
    .S1(net497),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_2 _42457_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(net489),
    .S1(net497),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _42458_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(net489),
    .S1(net497),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_1 _42459_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(net489),
    .S1(net497),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_2 _42460_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(net500),
    .S1(_00362_),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _42461_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(net489),
    .S1(net497),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_2 _42462_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(net489),
    .S1(net497),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_2 _42463_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(net489),
    .S1(net497),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_1 _42464_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(net489),
    .S1(net496),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_2 _42465_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(net489),
    .S1(net497),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_2 _42466_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(net500),
    .S1(_00362_),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_1 _42467_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(net478),
    .S1(net491),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_2 _42468_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(net480),
    .S1(net491),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_2 _42469_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(net481),
    .S1(net492),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_1 _42470_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(net480),
    .S1(net491),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _42471_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(net481),
    .S1(net491),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_2 _42472_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(net498),
    .S1(net502),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_2 _42473_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(net481),
    .S1(net491),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_2 _42474_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(net481),
    .S1(net491),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_2 _42475_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(net481),
    .S1(net492),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_1 _42476_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(net481),
    .S1(net491),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_2 _42477_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(net481),
    .S1(net491),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_2 _42478_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(net498),
    .S1(net502),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _42479_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(net478),
    .S1(net492),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_1 _42480_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(net481),
    .S1(net492),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_1 _42481_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(net481),
    .S1(net492),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_2 _42482_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(net481),
    .S1(net492),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_2 _42483_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(net481),
    .S1(net492),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_2 _42484_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(net498),
    .S1(net502),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_1 _42485_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(net478),
    .S1(net492),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_2 _42486_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(net481),
    .S1(net491),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_2 _42487_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(net481),
    .S1(net492),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_2 _42488_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(net481),
    .S1(net491),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _42489_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(net481),
    .S1(net492),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_2 _42490_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(net498),
    .S1(net502),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _42491_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(net478),
    .S1(net492),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_2 _42492_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(net488),
    .S1(net497),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_1 _42493_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(net488),
    .S1(net492),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_1 _42494_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(net488),
    .S1(net492),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_2 _42495_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(net488),
    .S1(net492),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_2 _42496_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(net500),
    .S1(net502),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _42497_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(net478),
    .S1(net492),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_2 _42498_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(net488),
    .S1(net497),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_2 _42499_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(net488),
    .S1(net492),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _42500_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(net488),
    .S1(net492),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_2 _42501_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(net488),
    .S1(net492),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_2 _42502_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(net500),
    .S1(net502),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_2 _42503_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(net486),
    .S1(net495),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_1 _42504_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(net486),
    .S1(net496),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_2 _42505_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(net486),
    .S1(net496),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_2 _42506_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(net486),
    .S1(net495),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_1 _42507_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(net486),
    .S1(net496),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_2 _42508_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(net499),
    .S1(net501),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_2 _42509_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(net486),
    .S1(net495),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_1 _42510_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(net485),
    .S1(net495),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_2 _42511_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(net485),
    .S1(net494),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_2 _42512_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(net483),
    .S1(net494),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _42513_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(net485),
    .S1(net495),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_2 _42514_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(net499),
    .S1(net501),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_2 _42515_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(net483),
    .S1(net494),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_2 _42516_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(net482),
    .S1(net494),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_2 _42517_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(net482),
    .S1(net494),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_2 _42518_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(net482),
    .S1(net494),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _42519_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(net482),
    .S1(net494),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_2 _42520_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(net499),
    .S1(net501),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_2 _42521_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(net483),
    .S1(net494),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_2 _42522_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(net482),
    .S1(net494),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_1 _42523_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(net482),
    .S1(net494),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_2 _42524_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(net482),
    .S1(net494),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_1 _42525_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(net482),
    .S1(net494),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_2 _42526_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(net499),
    .S1(net501),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_2 _42527_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(net483),
    .S1(net494),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_2 _42528_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(net482),
    .S1(net494),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_1 _42529_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(net482),
    .S1(net494),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_2 _42530_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(net482),
    .S1(net494),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_1 _42531_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(net482),
    .S1(net494),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_2 _42532_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(net499),
    .S1(net501),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_1 _42533_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(net486),
    .S1(net495),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_2 _42534_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(net485),
    .S1(net495),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_2 _42535_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(net485),
    .S1(net495),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_2 _42536_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(net486),
    .S1(net495),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _42537_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(net485),
    .S1(net495),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_2 _42538_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(net499),
    .S1(net501),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_2 _42539_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(net483),
    .S1(net493),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_2 _42540_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(net483),
    .S1(net493),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_1 _42541_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(net485),
    .S1(net493),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_2 _42542_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(net485),
    .S1(net493),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_2 _42543_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(net485),
    .S1(net493),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_2 _42544_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(net499),
    .S1(net501),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_2 _42545_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(net484),
    .S1(net495),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_1 _42546_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(net484),
    .S1(net493),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_2 _42547_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(net484),
    .S1(net493),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_1 _42548_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(net484),
    .S1(net493),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_2 _42549_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(net484),
    .S1(net493),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_2 _42550_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(net499),
    .S1(net501),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_2 _42551_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(net482),
    .S1(net494),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_2 _42552_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(net483),
    .S1(net493),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_1 _42553_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(net485),
    .S1(net493),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_2 _42554_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(net483),
    .S1(net493),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_2 _42555_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(net483),
    .S1(net493),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_2 _42556_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(net499),
    .S1(net501),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_2 _42557_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(net483),
    .S1(net494),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_2 _42558_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(net483),
    .S1(net493),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_1 _42559_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(net485),
    .S1(net493),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_2 _42560_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(net483),
    .S1(net493),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_2 _42561_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(net483),
    .S1(net494),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_2 _42562_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(net499),
    .S1(net501),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_2 _42563_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(net485),
    .S1(net495),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_1 _42564_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(net484),
    .S1(net493),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_2 _42565_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(net484),
    .S1(net493),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_1 _42566_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(net484),
    .S1(net493),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_2 _42567_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(net485),
    .S1(net493),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_2 _42568_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(net499),
    .S1(net501),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_2 _42569_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(net484),
    .S1(net495),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_2 _42570_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(net487),
    .S1(net495),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_2 _42571_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(net484),
    .S1(net495),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_1 _42572_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(net484),
    .S1(net495),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_2 _42573_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(net484),
    .S1(net495),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_2 _42574_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(net499),
    .S1(net501),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_2 _42575_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(net486),
    .S1(net496),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_1 _42576_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(net486),
    .S1(net496),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_2 _42577_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(net486),
    .S1(net496),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_2 _42578_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(net486),
    .S1(net496),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _42579_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(net486),
    .S1(net496),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_2 _42580_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(net500),
    .S1(net501),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _42581_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(net478),
    .S1(net491),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_2 _42582_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(net478),
    .S1(net492),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_2 _42583_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(net478),
    .S1(net492),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_1 _42584_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(net478),
    .S1(net492),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_2 _42585_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(net478),
    .S1(net491),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_2 _42586_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(net498),
    .S1(net502),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _42587_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(net436),
    .S1(net458),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _42588_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(net436),
    .S1(net458),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _42589_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(net436),
    .S1(net458),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _42590_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(net436),
    .S1(net458),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _42591_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(net436),
    .S1(net458),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _42592_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(net436),
    .S1(net458),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _42593_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(net436),
    .S1(net458),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _42594_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(net436),
    .S1(net458),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _42595_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(net436),
    .S1(net458),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _42596_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(net436),
    .S1(net458),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _42597_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(net436),
    .S1(net458),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _42598_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(net436),
    .S1(net458),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_2 _42599_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(net436),
    .S1(net458),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_2 _42600_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(net436),
    .S1(net458),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _42601_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(net436),
    .S1(net458),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _42602_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(net436),
    .S1(net458),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _42603_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(net436),
    .S1(net458),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _42604_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(_21107_),
    .S1(net458),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _42605_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(_21107_),
    .S1(net459),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _42606_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(_21107_),
    .S1(net459),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _42607_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_21107_),
    .S1(net459),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _42608_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_21107_),
    .S1(net459),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _42609_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_21107_),
    .S1(net459),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _42610_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_21107_),
    .S1(net459),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _42611_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_21107_),
    .S1(net459),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _42612_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_21107_),
    .S1(net459),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _42613_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_21107_),
    .S1(net459),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _42614_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_21107_),
    .S1(net459),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _42615_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_21107_),
    .S1(net459),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_1 _42616_ (.D(_02687_),
    .Q(\alu_shl[0] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 _42617_ (.D(_02688_),
    .Q(\alu_shl[1] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42618_ (.D(_02689_),
    .Q(\alu_shl[2] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 _42619_ (.D(_02690_),
    .Q(\alu_shl[3] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 _42620_ (.D(_02691_),
    .Q(\alu_shl[4] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42621_ (.D(_02692_),
    .Q(\alu_shl[5] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42622_ (.D(_02693_),
    .Q(\alu_shl[6] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42623_ (.D(_02694_),
    .Q(\alu_shl[7] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42624_ (.D(_02695_),
    .Q(\alu_shl[8] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42625_ (.D(_02696_),
    .Q(\alu_shl[9] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42626_ (.D(_02697_),
    .Q(\alu_shl[10] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42627_ (.D(_02698_),
    .Q(\alu_shl[11] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 _42628_ (.D(_02699_),
    .Q(\alu_shl[12] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42629_ (.D(_02700_),
    .Q(\alu_shl[13] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42630_ (.D(_02701_),
    .Q(\alu_shl[14] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42631_ (.D(_02702_),
    .Q(\alu_shl[15] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _42632_ (.D(_02703_),
    .Q(alu_wait),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _42633_ (.D(_02704_),
    .Q(\latched_rd[3] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _42634_ (.D(_02705_),
    .Q(\latched_rd[2] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42635_ (.D(_02706_),
    .Q(\latched_rd[1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42636_ (.D(_02707_),
    .Q(\latched_rd[0] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_4 _42637_ (.D(_02708_),
    .Q(\decoded_imm[31] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_4 _42638_ (.D(_02709_),
    .Q(\decoded_imm[30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _42639_ (.D(_02710_),
    .Q(\decoded_imm[29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42640_ (.D(_02711_),
    .Q(\decoded_imm[28] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_4 _42641_ (.D(_02712_),
    .Q(\decoded_imm[27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_4 _42642_ (.D(_02713_),
    .Q(\decoded_imm[26] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42643_ (.D(_02714_),
    .Q(\decoded_imm[25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42644_ (.D(_02715_),
    .Q(\decoded_imm[24] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42645_ (.D(_02716_),
    .Q(\decoded_imm[23] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42646_ (.D(_02717_),
    .Q(\decoded_imm[22] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42647_ (.D(_02718_),
    .Q(\decoded_imm[21] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42648_ (.D(_02719_),
    .Q(\decoded_imm[20] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42649_ (.D(_02720_),
    .Q(\decoded_imm[19] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _42650_ (.D(_02721_),
    .Q(\decoded_imm[18] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _42651_ (.D(_02722_),
    .Q(\decoded_imm[17] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_2 _42652_ (.D(_02723_),
    .Q(\decoded_imm[16] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_2 _42653_ (.D(_02724_),
    .Q(\decoded_imm[15] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _42654_ (.D(_02725_),
    .Q(\decoded_imm[14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42655_ (.D(_02726_),
    .Q(\decoded_imm[13] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_4 _42656_ (.D(_02727_),
    .Q(\decoded_imm[12] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42657_ (.D(_02728_),
    .Q(\decoded_imm[11] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42658_ (.D(_02729_),
    .Q(\decoded_imm[10] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_2 _42659_ (.D(_02730_),
    .Q(\decoded_imm[9] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42660_ (.D(_02731_),
    .Q(\decoded_imm[8] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42661_ (.D(_02732_),
    .Q(\decoded_imm[7] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_2 _42662_ (.D(_02733_),
    .Q(\decoded_imm[6] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_2 _42663_ (.D(_02734_),
    .Q(\decoded_imm[5] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 _42664_ (.D(_02735_),
    .Q(\decoded_imm[4] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42665_ (.D(_02736_),
    .Q(\decoded_imm[3] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _42666_ (.D(_02737_),
    .Q(\decoded_imm[2] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42667_ (.D(_02738_),
    .Q(\decoded_imm[1] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _42668_ (.D(_02739_),
    .Q(\irq_pending[31] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _42669_ (.D(_02740_),
    .Q(\irq_pending[30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42670_ (.D(_02741_),
    .Q(\irq_pending[29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _42671_ (.D(_02742_),
    .Q(\irq_pending[28] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _42672_ (.D(_02743_),
    .Q(\irq_pending[27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _42673_ (.D(_02744_),
    .Q(\irq_pending[26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42674_ (.D(_02745_),
    .Q(\irq_pending[25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42675_ (.D(_02746_),
    .Q(\irq_pending[24] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _42676_ (.D(_02747_),
    .Q(\irq_pending[23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _42677_ (.D(_02748_),
    .Q(\irq_pending[22] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 _42678_ (.D(_02749_),
    .Q(\irq_pending[21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_2 _42679_ (.D(_02750_),
    .Q(\irq_pending[20] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42680_ (.D(_02751_),
    .Q(\irq_pending[19] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42681_ (.D(_02752_),
    .Q(\irq_pending[18] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42682_ (.D(_02753_),
    .Q(\irq_pending[17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _42683_ (.D(_02754_),
    .Q(\irq_pending[16] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _42684_ (.D(_02755_),
    .Q(\irq_pending[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42685_ (.D(_02756_),
    .Q(\irq_pending[14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42686_ (.D(_02757_),
    .Q(\irq_pending[13] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42687_ (.D(_02758_),
    .Q(\irq_pending[12] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _42688_ (.D(_02759_),
    .Q(\irq_pending[11] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _42689_ (.D(_02760_),
    .Q(\irq_pending[10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42690_ (.D(_02761_),
    .Q(\irq_pending[9] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42691_ (.D(_02762_),
    .Q(\irq_pending[8] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _42692_ (.D(_02763_),
    .Q(\irq_pending[7] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _42693_ (.D(_02764_),
    .Q(\irq_pending[6] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _42694_ (.D(_02765_),
    .Q(\irq_pending[5] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42695_ (.D(_02766_),
    .Q(\irq_pending[4] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42696_ (.D(_02767_),
    .Q(\irq_pending[3] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _42697_ (.D(_02768_),
    .Q(\irq_pending[1] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _42698_ (.D(_02769_),
    .Q(\irq_pending[0] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42699_ (.D(_02770_),
    .Q(\reg_next_pc[0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _42700_ (.D(_00045_),
    .Q(\mem_wordsize[0] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_2 _42701_ (.D(_00046_),
    .Q(\mem_wordsize[1] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _42702_ (.D(_00047_),
    .Q(\mem_wordsize[2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 _42703_ (.D(_21109_),
    .Q(\reg_out[0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _42704_ (.D(_21120_),
    .Q(\reg_out[1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _42705_ (.D(_21131_),
    .Q(\reg_out[2] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 _42706_ (.D(_21134_),
    .Q(\reg_out[3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _42707_ (.D(_21135_),
    .Q(\reg_out[4] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _42708_ (.D(_21136_),
    .Q(\reg_out[5] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _42709_ (.D(_21137_),
    .Q(\reg_out[6] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _42710_ (.D(_21138_),
    .Q(\reg_out[7] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _42711_ (.D(_21139_),
    .Q(\reg_out[8] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _42712_ (.D(_21140_),
    .Q(\reg_out[9] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _42713_ (.D(_21110_),
    .Q(\reg_out[10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _42714_ (.D(_21111_),
    .Q(\reg_out[11] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42715_ (.D(_21112_),
    .Q(\reg_out[12] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _42716_ (.D(_21113_),
    .Q(\reg_out[13] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_1 _42717_ (.D(_21114_),
    .Q(\reg_out[14] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _42718_ (.D(_21115_),
    .Q(\reg_out[15] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _42719_ (.D(_21116_),
    .Q(\reg_out[16] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_1 _42720_ (.D(_21117_),
    .Q(\reg_out[17] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _42721_ (.D(_21118_),
    .Q(\reg_out[18] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _42722_ (.D(_21119_),
    .Q(\reg_out[19] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_1 _42723_ (.D(_21121_),
    .Q(\reg_out[20] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_1 _42724_ (.D(_21122_),
    .Q(\reg_out[21] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _42725_ (.D(_21123_),
    .Q(\reg_out[22] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _42726_ (.D(_21124_),
    .Q(\reg_out[23] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _42727_ (.D(_21125_),
    .Q(\reg_out[24] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _42728_ (.D(_21126_),
    .Q(\reg_out[25] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _42729_ (.D(_21127_),
    .Q(\reg_out[26] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _42730_ (.D(_21128_),
    .Q(\reg_out[27] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _42731_ (.D(_21129_),
    .Q(\reg_out[28] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _42732_ (.D(_21130_),
    .Q(\reg_out[29] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42733_ (.D(_21132_),
    .Q(\reg_out[30] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _42734_ (.D(_21133_),
    .Q(\reg_out[31] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _42735_ (.D(_00004_),
    .Q(\irq_pending[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42736_ (.D(_00003_),
    .Q(decoder_trigger),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _42737_ (.D(\alu_out[0] ),
    .Q(\alu_out_q[0] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 _42738_ (.D(\alu_out[1] ),
    .Q(\alu_out_q[1] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42739_ (.D(\alu_out[2] ),
    .Q(\alu_out_q[2] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42740_ (.D(\alu_out[3] ),
    .Q(\alu_out_q[3] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42741_ (.D(\alu_out[4] ),
    .Q(\alu_out_q[4] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 _42742_ (.D(\alu_out[5] ),
    .Q(\alu_out_q[5] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 _42743_ (.D(\alu_out[6] ),
    .Q(\alu_out_q[6] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 _42744_ (.D(\alu_out[7] ),
    .Q(\alu_out_q[7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 _42745_ (.D(\alu_out[8] ),
    .Q(\alu_out_q[8] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 _42746_ (.D(\alu_out[9] ),
    .Q(\alu_out_q[9] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42747_ (.D(\alu_out[10] ),
    .Q(\alu_out_q[10] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42748_ (.D(\alu_out[11] ),
    .Q(\alu_out_q[11] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42749_ (.D(\alu_out[12] ),
    .Q(\alu_out_q[12] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 _42750_ (.D(\alu_out[13] ),
    .Q(\alu_out_q[13] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 _42751_ (.D(\alu_out[14] ),
    .Q(\alu_out_q[14] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42752_ (.D(\alu_out[15] ),
    .Q(\alu_out_q[15] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42753_ (.D(\alu_out[16] ),
    .Q(\alu_out_q[16] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42754_ (.D(\alu_out[17] ),
    .Q(\alu_out_q[17] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42755_ (.D(\alu_out[18] ),
    .Q(\alu_out_q[18] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42756_ (.D(\alu_out[19] ),
    .Q(\alu_out_q[19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42757_ (.D(\alu_out[20] ),
    .Q(\alu_out_q[20] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42758_ (.D(\alu_out[21] ),
    .Q(\alu_out_q[21] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42759_ (.D(\alu_out[22] ),
    .Q(\alu_out_q[22] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42760_ (.D(\alu_out[23] ),
    .Q(\alu_out_q[23] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42761_ (.D(\alu_out[24] ),
    .Q(\alu_out_q[24] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42762_ (.D(\alu_out[25] ),
    .Q(\alu_out_q[25] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42763_ (.D(\alu_out[26] ),
    .Q(\alu_out_q[26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42764_ (.D(\alu_out[27] ),
    .Q(\alu_out_q[27] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_2 _42765_ (.D(\alu_out[28] ),
    .Q(\alu_out_q[28] ),
    .CLK(clknet_5_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42766_ (.D(\alu_out[29] ),
    .Q(\alu_out_q[29] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _42767_ (.D(\alu_out[30] ),
    .Q(\alu_out_q[30] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _42768_ (.D(\alu_out[31] ),
    .Q(\alu_out_q[31] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_4 _42769_ (.D(_00005_),
    .Q(is_lui_auipc_jal),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _42770_ (.D(_00006_),
    .Q(is_slti_blt_slt),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _42771_ (.D(_00007_),
    .Q(is_sltiu_bltu_sltu),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _42772_ (.D(_02591_),
    .Q(\alu_add_sub[0] ),
    .CLK(clknet_5_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42773_ (.D(_02602_),
    .Q(\alu_add_sub[1] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 _42774_ (.D(_02613_),
    .Q(\alu_add_sub[2] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 _42775_ (.D(_02616_),
    .Q(\alu_add_sub[3] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42776_ (.D(_02617_),
    .Q(\alu_add_sub[4] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42777_ (.D(_02618_),
    .Q(\alu_add_sub[5] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 _42778_ (.D(_02619_),
    .Q(\alu_add_sub[6] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 _42779_ (.D(_02620_),
    .Q(\alu_add_sub[7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 _42780_ (.D(_02621_),
    .Q(\alu_add_sub[8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42781_ (.D(_02622_),
    .Q(\alu_add_sub[9] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42782_ (.D(_02592_),
    .Q(\alu_add_sub[10] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42783_ (.D(_02593_),
    .Q(\alu_add_sub[11] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42784_ (.D(_02594_),
    .Q(\alu_add_sub[12] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _42785_ (.D(_02595_),
    .Q(\alu_add_sub[13] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 _42786_ (.D(_02596_),
    .Q(\alu_add_sub[14] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 _42787_ (.D(_02597_),
    .Q(\alu_add_sub[15] ),
    .CLK(clknet_5_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42788_ (.D(_02598_),
    .Q(\alu_add_sub[16] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42789_ (.D(_02599_),
    .Q(\alu_add_sub[17] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42790_ (.D(_02600_),
    .Q(\alu_add_sub[18] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42791_ (.D(_02601_),
    .Q(\alu_add_sub[19] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _42792_ (.D(_02603_),
    .Q(\alu_add_sub[20] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _42793_ (.D(_02604_),
    .Q(\alu_add_sub[21] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _42794_ (.D(_02605_),
    .Q(\alu_add_sub[22] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42795_ (.D(_02606_),
    .Q(\alu_add_sub[23] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42796_ (.D(_02607_),
    .Q(\alu_add_sub[24] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42797_ (.D(_02608_),
    .Q(\alu_add_sub[25] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42798_ (.D(_02609_),
    .Q(\alu_add_sub[26] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _42799_ (.D(_02610_),
    .Q(\alu_add_sub[27] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _42800_ (.D(_02611_),
    .Q(\alu_add_sub[28] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _42801_ (.D(_02612_),
    .Q(\alu_add_sub[29] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _42802_ (.D(_02614_),
    .Q(\alu_add_sub[30] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _42803_ (.D(_02615_),
    .Q(\alu_add_sub[31] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _42804_ (.D(_21144_),
    .Q(\alu_shl[16] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 _42805_ (.D(_21145_),
    .Q(\alu_shl[17] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42806_ (.D(_21146_),
    .Q(\alu_shl[18] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42807_ (.D(_21147_),
    .Q(\alu_shl[19] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42808_ (.D(_21148_),
    .Q(\alu_shl[20] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42809_ (.D(_21149_),
    .Q(\alu_shl[21] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42810_ (.D(_21150_),
    .Q(\alu_shl[22] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42811_ (.D(_21151_),
    .Q(\alu_shl[23] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42812_ (.D(_21152_),
    .Q(\alu_shl[24] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42813_ (.D(_21153_),
    .Q(\alu_shl[25] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42814_ (.D(_21154_),
    .Q(\alu_shl[26] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42815_ (.D(_21155_),
    .Q(\alu_shl[27] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42816_ (.D(_21156_),
    .Q(\alu_shl[28] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42817_ (.D(_21157_),
    .Q(\alu_shl[29] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42818_ (.D(_21158_),
    .Q(\alu_shl[30] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42819_ (.D(_21159_),
    .Q(\alu_shl[31] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42820_ (.D(_21160_),
    .Q(\alu_shr[0] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 _42821_ (.D(_21171_),
    .Q(\alu_shr[1] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42822_ (.D(_21182_),
    .Q(\alu_shr[2] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42823_ (.D(_21185_),
    .Q(\alu_shr[3] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42824_ (.D(_21186_),
    .Q(\alu_shr[4] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 _42825_ (.D(_21187_),
    .Q(\alu_shr[5] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42826_ (.D(_21188_),
    .Q(\alu_shr[6] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _42827_ (.D(_21189_),
    .Q(\alu_shr[7] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42828_ (.D(_21190_),
    .Q(\alu_shr[8] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42829_ (.D(_21191_),
    .Q(\alu_shr[9] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42830_ (.D(_21161_),
    .Q(\alu_shr[10] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42831_ (.D(_21162_),
    .Q(\alu_shr[11] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _42832_ (.D(_21163_),
    .Q(\alu_shr[12] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42833_ (.D(_21164_),
    .Q(\alu_shr[13] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42834_ (.D(_21165_),
    .Q(\alu_shr[14] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42835_ (.D(_21166_),
    .Q(\alu_shr[15] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _42836_ (.D(_21167_),
    .Q(\alu_shr[16] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42837_ (.D(_21168_),
    .Q(\alu_shr[17] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42838_ (.D(_21169_),
    .Q(\alu_shr[18] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42839_ (.D(_21170_),
    .Q(\alu_shr[19] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42840_ (.D(_21172_),
    .Q(\alu_shr[20] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42841_ (.D(_21173_),
    .Q(\alu_shr[21] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42842_ (.D(_21174_),
    .Q(\alu_shr[22] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42843_ (.D(_21175_),
    .Q(\alu_shr[23] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42844_ (.D(_21176_),
    .Q(\alu_shr[24] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42845_ (.D(_21177_),
    .Q(\alu_shr[25] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42846_ (.D(_21178_),
    .Q(\alu_shr[26] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42847_ (.D(_21179_),
    .Q(\alu_shr[27] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42848_ (.D(_21180_),
    .Q(\alu_shr[28] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42849_ (.D(_21181_),
    .Q(\alu_shr[29] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42850_ (.D(_21183_),
    .Q(\alu_shr[30] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _42851_ (.D(_21184_),
    .Q(\alu_shr[31] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42852_ (.D(_00000_),
    .Q(alu_eq),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42853_ (.D(_00002_),
    .Q(alu_ltu),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42854_ (.D(_00001_),
    .Q(alu_lts),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 _42855_ (.D(_02623_),
    .Q(\pcpi_mul.rd[0] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 _42856_ (.D(_02624_),
    .Q(\pcpi_mul.rd[1] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 _42857_ (.D(_02625_),
    .Q(\pcpi_mul.rd[2] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _42858_ (.D(_02626_),
    .Q(\pcpi_mul.rd[3] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _42859_ (.D(_02627_),
    .Q(\pcpi_mul.rd[4] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 _42860_ (.D(_02628_),
    .Q(\pcpi_mul.rd[5] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 _42861_ (.D(_02683_),
    .Q(\pcpi_mul.rd[6] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _42862_ (.D(_02684_),
    .Q(\pcpi_mul.rd[7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _42863_ (.D(_02685_),
    .Q(\pcpi_mul.rd[8] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42864_ (.D(_02686_),
    .Q(\pcpi_mul.rd[9] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42865_ (.D(_02629_),
    .Q(\pcpi_mul.rd[10] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _42866_ (.D(_02630_),
    .Q(\pcpi_mul.rd[11] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42867_ (.D(_02631_),
    .Q(\pcpi_mul.rd[12] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42868_ (.D(_02632_),
    .Q(\pcpi_mul.rd[13] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42869_ (.D(_02633_),
    .Q(\pcpi_mul.rd[14] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42870_ (.D(_02634_),
    .Q(\pcpi_mul.rd[15] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_4 _42871_ (.D(_02635_),
    .Q(\pcpi_mul.rd[16] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_4 _42872_ (.D(_02636_),
    .Q(\pcpi_mul.rd[17] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_4 _42873_ (.D(_02637_),
    .Q(\pcpi_mul.rd[18] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_4 _42874_ (.D(_02638_),
    .Q(\pcpi_mul.rd[19] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_4 _42875_ (.D(_02639_),
    .Q(\pcpi_mul.rd[20] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_4 _42876_ (.D(_02640_),
    .Q(\pcpi_mul.rd[21] ),
    .CLK(clknet_5_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _42877_ (.D(_02641_),
    .Q(\pcpi_mul.rd[22] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_4 _42878_ (.D(_02642_),
    .Q(\pcpi_mul.rd[23] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _42879_ (.D(_02643_),
    .Q(\pcpi_mul.rd[24] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 _42880_ (.D(_02644_),
    .Q(\pcpi_mul.rd[25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_1 _42881_ (.D(_02645_),
    .Q(\pcpi_mul.rd[26] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42882_ (.D(_02646_),
    .Q(\pcpi_mul.rd[27] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42883_ (.D(_02647_),
    .Q(\pcpi_mul.rd[28] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 _42884_ (.D(_02648_),
    .Q(\pcpi_mul.rd[29] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 _42885_ (.D(_02649_),
    .Q(\pcpi_mul.rd[30] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 _42886_ (.D(_02650_),
    .Q(\pcpi_mul.rd[31] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 _42887_ (.D(_02651_),
    .Q(\pcpi_mul.rd[32] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 _42888_ (.D(_02652_),
    .Q(\pcpi_mul.rd[33] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 _42889_ (.D(_02653_),
    .Q(\pcpi_mul.rd[34] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _42890_ (.D(_02654_),
    .Q(\pcpi_mul.rd[35] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _42891_ (.D(_02655_),
    .Q(\pcpi_mul.rd[36] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42892_ (.D(_02656_),
    .Q(\pcpi_mul.rd[37] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42893_ (.D(_02657_),
    .Q(\pcpi_mul.rd[38] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42894_ (.D(_02658_),
    .Q(\pcpi_mul.rd[39] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _42895_ (.D(_02659_),
    .Q(\pcpi_mul.rd[40] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _42896_ (.D(_02660_),
    .Q(\pcpi_mul.rd[41] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42897_ (.D(_02661_),
    .Q(\pcpi_mul.rd[42] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42898_ (.D(_02662_),
    .Q(\pcpi_mul.rd[43] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _42899_ (.D(_02663_),
    .Q(\pcpi_mul.rd[44] ),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42900_ (.D(_02664_),
    .Q(\pcpi_mul.rd[45] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _42901_ (.D(_02665_),
    .Q(\pcpi_mul.rd[46] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_4 _42902_ (.D(_02666_),
    .Q(\pcpi_mul.rd[47] ),
    .CLK(clknet_opt_10_clk));
 sky130_fd_sc_hd__dfxtp_4 _42903_ (.D(_02667_),
    .Q(\pcpi_mul.rd[48] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_4 _42904_ (.D(_02668_),
    .Q(\pcpi_mul.rd[49] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_4 _42905_ (.D(_02669_),
    .Q(\pcpi_mul.rd[50] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_4 _42906_ (.D(_02670_),
    .Q(\pcpi_mul.rd[51] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 _42907_ (.D(_02671_),
    .Q(\pcpi_mul.rd[52] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 _42908_ (.D(_02672_),
    .Q(\pcpi_mul.rd[53] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 _42909_ (.D(_02673_),
    .Q(\pcpi_mul.rd[54] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _42910_ (.D(_02674_),
    .Q(\pcpi_mul.rd[55] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _42911_ (.D(_02675_),
    .Q(\pcpi_mul.rd[56] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_4 _42912_ (.D(_02676_),
    .Q(\pcpi_mul.rd[57] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _42913_ (.D(_02677_),
    .Q(\pcpi_mul.rd[58] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42914_ (.D(_02678_),
    .Q(\pcpi_mul.rd[59] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42915_ (.D(_02679_),
    .Q(\pcpi_mul.rd[60] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 _42916_ (.D(_02680_),
    .Q(\pcpi_mul.rd[61] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42917_ (.D(_02681_),
    .Q(\pcpi_mul.rd[62] ),
    .CLK(clknet_5_23_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42918_ (.D(_02682_),
    .Q(\pcpi_mul.rd[63] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_4 _42919_ (.D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 _42920_ (.D(_00038_),
    .Q(\cpu_state[0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _42921_ (.D(_00039_),
    .Q(\cpu_state[1] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _42922_ (.D(_00040_),
    .Q(\cpu_state[2] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_4 _42923_ (.D(_00041_),
    .Q(\cpu_state[3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_4 _42924_ (.D(_00042_),
    .Q(\cpu_state[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_4 _42925_ (.D(_00043_),
    .Q(\cpu_state[5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _42926_ (.D(_00044_),
    .Q(\cpu_state[6] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42927_ (.D(_02771_),
    .Q(\cpuregs[8][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _42928_ (.D(_02772_),
    .Q(\cpuregs[8][1] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _42929_ (.D(_02773_),
    .Q(\cpuregs[8][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _42930_ (.D(_02774_),
    .Q(\cpuregs[8][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42931_ (.D(_02775_),
    .Q(\cpuregs[8][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _42932_ (.D(_02776_),
    .Q(\cpuregs[8][5] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42933_ (.D(_02777_),
    .Q(\cpuregs[8][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42934_ (.D(_02778_),
    .Q(\cpuregs[8][7] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42935_ (.D(_02779_),
    .Q(\cpuregs[8][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _42936_ (.D(_02780_),
    .Q(\cpuregs[8][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _42937_ (.D(_02781_),
    .Q(\cpuregs[8][10] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _42938_ (.D(_02782_),
    .Q(\cpuregs[8][11] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _42939_ (.D(_02783_),
    .Q(\cpuregs[8][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42940_ (.D(_02784_),
    .Q(\cpuregs[8][13] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _42941_ (.D(_02785_),
    .Q(\cpuregs[8][14] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _42942_ (.D(_02786_),
    .Q(\cpuregs[8][15] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _42943_ (.D(_02787_),
    .Q(\cpuregs[8][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42944_ (.D(_02788_),
    .Q(\cpuregs[8][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _42945_ (.D(_02789_),
    .Q(\cpuregs[8][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _42946_ (.D(_02790_),
    .Q(\cpuregs[8][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _42947_ (.D(_02791_),
    .Q(\cpuregs[8][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _42948_ (.D(_02792_),
    .Q(\cpuregs[8][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _42949_ (.D(_02793_),
    .Q(\cpuregs[8][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _42950_ (.D(_02794_),
    .Q(\cpuregs[8][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42951_ (.D(_02795_),
    .Q(\cpuregs[8][24] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _42952_ (.D(_02796_),
    .Q(\cpuregs[8][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _42953_ (.D(_02797_),
    .Q(\cpuregs[8][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42954_ (.D(_02798_),
    .Q(\cpuregs[8][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _42955_ (.D(_02799_),
    .Q(\cpuregs[8][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _42956_ (.D(_02800_),
    .Q(\cpuregs[8][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _42957_ (.D(_02801_),
    .Q(\cpuregs[8][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _42958_ (.D(_02802_),
    .Q(\cpuregs[8][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _42959_ (.D(_02803_),
    .Q(\cpuregs[14][0] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _42960_ (.D(_02804_),
    .Q(\cpuregs[14][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42961_ (.D(_02805_),
    .Q(\cpuregs[14][2] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42962_ (.D(_02806_),
    .Q(\cpuregs[14][3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _42963_ (.D(_02807_),
    .Q(\cpuregs[14][4] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _42964_ (.D(_02808_),
    .Q(\cpuregs[14][5] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _42965_ (.D(_02809_),
    .Q(\cpuregs[14][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42966_ (.D(_02810_),
    .Q(\cpuregs[14][7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _42967_ (.D(_02811_),
    .Q(\cpuregs[14][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _42968_ (.D(_02812_),
    .Q(\cpuregs[14][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _42969_ (.D(_02813_),
    .Q(\cpuregs[14][10] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _42970_ (.D(_02814_),
    .Q(\cpuregs[14][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _42971_ (.D(_02815_),
    .Q(\cpuregs[14][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42972_ (.D(_02816_),
    .Q(\cpuregs[14][13] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _42973_ (.D(_02817_),
    .Q(\cpuregs[14][14] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _42974_ (.D(_02818_),
    .Q(\cpuregs[14][15] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42975_ (.D(_02819_),
    .Q(\cpuregs[14][16] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _42976_ (.D(_02820_),
    .Q(\cpuregs[14][17] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _42977_ (.D(_02821_),
    .Q(\cpuregs[14][18] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _42978_ (.D(_02822_),
    .Q(\cpuregs[14][19] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _42979_ (.D(_02823_),
    .Q(\cpuregs[14][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _42980_ (.D(_02824_),
    .Q(\cpuregs[14][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _42981_ (.D(_02825_),
    .Q(\cpuregs[14][22] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _42982_ (.D(_02826_),
    .Q(\cpuregs[14][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42983_ (.D(_02827_),
    .Q(\cpuregs[14][24] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42984_ (.D(_02828_),
    .Q(\cpuregs[14][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _42985_ (.D(_02829_),
    .Q(\cpuregs[14][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _42986_ (.D(_02830_),
    .Q(\cpuregs[14][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _42987_ (.D(_02831_),
    .Q(\cpuregs[14][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _42988_ (.D(_02832_),
    .Q(\cpuregs[14][29] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _42989_ (.D(_02833_),
    .Q(\cpuregs[14][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _42990_ (.D(_02834_),
    .Q(\cpuregs[14][31] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _42991_ (.D(_02835_),
    .Q(\cpuregs[0][0] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _42992_ (.D(_02836_),
    .Q(\cpuregs[0][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42993_ (.D(_02837_),
    .Q(\cpuregs[0][2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42994_ (.D(_02838_),
    .Q(\cpuregs[0][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42995_ (.D(_02839_),
    .Q(\cpuregs[0][4] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _42996_ (.D(_02840_),
    .Q(\cpuregs[0][5] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _42997_ (.D(_02841_),
    .Q(\cpuregs[0][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42998_ (.D(_02842_),
    .Q(\cpuregs[0][7] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _42999_ (.D(_02843_),
    .Q(\cpuregs[0][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43000_ (.D(_02844_),
    .Q(\cpuregs[0][9] ),
    .CLK(clknet_5_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43001_ (.D(_02845_),
    .Q(\cpuregs[0][10] ),
    .CLK(clknet_5_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43002_ (.D(_02846_),
    .Q(\cpuregs[0][11] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43003_ (.D(_02847_),
    .Q(\cpuregs[0][12] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43004_ (.D(_02848_),
    .Q(\cpuregs[0][13] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _43005_ (.D(_02849_),
    .Q(\cpuregs[0][14] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43006_ (.D(_02850_),
    .Q(\cpuregs[0][15] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43007_ (.D(_02851_),
    .Q(\cpuregs[0][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43008_ (.D(_02852_),
    .Q(\cpuregs[0][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43009_ (.D(_02853_),
    .Q(\cpuregs[0][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43010_ (.D(_02854_),
    .Q(\cpuregs[0][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43011_ (.D(_02855_),
    .Q(\cpuregs[0][20] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43012_ (.D(_02856_),
    .Q(\cpuregs[0][21] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_1 _43013_ (.D(_02857_),
    .Q(\cpuregs[0][22] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43014_ (.D(_02858_),
    .Q(\cpuregs[0][23] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43015_ (.D(_02859_),
    .Q(\cpuregs[0][24] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _43016_ (.D(_02860_),
    .Q(\cpuregs[0][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43017_ (.D(_02861_),
    .Q(\cpuregs[0][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43018_ (.D(_02862_),
    .Q(\cpuregs[0][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43019_ (.D(_02863_),
    .Q(\cpuregs[0][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43020_ (.D(_02864_),
    .Q(\cpuregs[0][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43021_ (.D(_02865_),
    .Q(\cpuregs[0][30] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43022_ (.D(_02866_),
    .Q(\cpuregs[0][31] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43023_ (.D(_02867_),
    .Q(\cpuregs[10][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43024_ (.D(_02868_),
    .Q(\cpuregs[10][1] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _43025_ (.D(_02869_),
    .Q(\cpuregs[10][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43026_ (.D(_02870_),
    .Q(\cpuregs[10][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43027_ (.D(_02871_),
    .Q(\cpuregs[10][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43028_ (.D(_02872_),
    .Q(\cpuregs[10][5] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43029_ (.D(_02873_),
    .Q(\cpuregs[10][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43030_ (.D(_02874_),
    .Q(\cpuregs[10][7] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43031_ (.D(_02875_),
    .Q(\cpuregs[10][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43032_ (.D(_02876_),
    .Q(\cpuregs[10][9] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43033_ (.D(_02877_),
    .Q(\cpuregs[10][10] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43034_ (.D(_02878_),
    .Q(\cpuregs[10][11] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43035_ (.D(_02879_),
    .Q(\cpuregs[10][12] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43036_ (.D(_02880_),
    .Q(\cpuregs[10][13] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43037_ (.D(_02881_),
    .Q(\cpuregs[10][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43038_ (.D(_02882_),
    .Q(\cpuregs[10][15] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43039_ (.D(_02883_),
    .Q(\cpuregs[10][16] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _43040_ (.D(_02884_),
    .Q(\cpuregs[10][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43041_ (.D(_02885_),
    .Q(\cpuregs[10][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43042_ (.D(_02886_),
    .Q(\cpuregs[10][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43043_ (.D(_02887_),
    .Q(\cpuregs[10][20] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43044_ (.D(_02888_),
    .Q(\cpuregs[10][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43045_ (.D(_02889_),
    .Q(\cpuregs[10][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43046_ (.D(_02890_),
    .Q(\cpuregs[10][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43047_ (.D(_02891_),
    .Q(\cpuregs[10][24] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _43048_ (.D(_02892_),
    .Q(\cpuregs[10][25] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43049_ (.D(_02893_),
    .Q(\cpuregs[10][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43050_ (.D(_02894_),
    .Q(\cpuregs[10][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43051_ (.D(_02895_),
    .Q(\cpuregs[10][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43052_ (.D(_02896_),
    .Q(\cpuregs[10][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43053_ (.D(_02897_),
    .Q(\cpuregs[10][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43054_ (.D(_02898_),
    .Q(\cpuregs[10][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43055_ (.D(_02899_),
    .Q(\cpuregs[18][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43056_ (.D(_02900_),
    .Q(\cpuregs[18][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43057_ (.D(_02901_),
    .Q(\cpuregs[18][2] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43058_ (.D(_02902_),
    .Q(\cpuregs[18][3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43059_ (.D(_02903_),
    .Q(\cpuregs[18][4] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43060_ (.D(_02904_),
    .Q(\cpuregs[18][5] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43061_ (.D(_02905_),
    .Q(\cpuregs[18][6] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43062_ (.D(_02906_),
    .Q(\cpuregs[18][7] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43063_ (.D(_02907_),
    .Q(\cpuregs[18][8] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43064_ (.D(_02908_),
    .Q(\cpuregs[18][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43065_ (.D(_02909_),
    .Q(\cpuregs[18][10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43066_ (.D(_02910_),
    .Q(\cpuregs[18][11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43067_ (.D(_02911_),
    .Q(\cpuregs[18][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43068_ (.D(_02912_),
    .Q(\cpuregs[18][13] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43069_ (.D(_02913_),
    .Q(\cpuregs[18][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43070_ (.D(_02914_),
    .Q(\cpuregs[18][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43071_ (.D(_02915_),
    .Q(\cpuregs[18][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43072_ (.D(_02916_),
    .Q(\cpuregs[18][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43073_ (.D(_02917_),
    .Q(\cpuregs[18][18] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43074_ (.D(_02918_),
    .Q(\cpuregs[18][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43075_ (.D(_02919_),
    .Q(\cpuregs[18][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43076_ (.D(_02920_),
    .Q(\cpuregs[18][21] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43077_ (.D(_02921_),
    .Q(\cpuregs[18][22] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _43078_ (.D(_02922_),
    .Q(\cpuregs[18][23] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43079_ (.D(_02923_),
    .Q(\cpuregs[18][24] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _43080_ (.D(_02924_),
    .Q(\cpuregs[18][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43081_ (.D(_02925_),
    .Q(\cpuregs[18][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43082_ (.D(_02926_),
    .Q(\cpuregs[18][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43083_ (.D(_02927_),
    .Q(\cpuregs[18][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43084_ (.D(_02928_),
    .Q(\cpuregs[18][29] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43085_ (.D(_02929_),
    .Q(\cpuregs[18][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43086_ (.D(_02930_),
    .Q(\cpuregs[18][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43087_ (.D(_02931_),
    .Q(\mem_rdata_q[0] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _43088_ (.D(_02932_),
    .Q(\mem_rdata_q[1] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _43089_ (.D(_02933_),
    .Q(\mem_rdata_q[2] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _43090_ (.D(_02934_),
    .Q(\mem_rdata_q[3] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _43091_ (.D(_02935_),
    .Q(\mem_rdata_q[4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43092_ (.D(_02936_),
    .Q(\mem_rdata_q[5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 _43093_ (.D(_02937_),
    .Q(\mem_rdata_q[6] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_2 _43094_ (.D(_02938_),
    .Q(\mem_rdata_q[7] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _43095_ (.D(_02939_),
    .Q(\mem_rdata_q[8] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _43096_ (.D(_02940_),
    .Q(\mem_rdata_q[9] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43097_ (.D(_02941_),
    .Q(\mem_rdata_q[10] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _43098_ (.D(_02942_),
    .Q(\mem_rdata_q[11] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _43099_ (.D(_02943_),
    .Q(\mem_rdata_q[12] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _43100_ (.D(_02944_),
    .Q(\mem_rdata_q[13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 _43101_ (.D(_02945_),
    .Q(\mem_rdata_q[14] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _43102_ (.D(_02946_),
    .Q(\mem_rdata_q[15] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 _43103_ (.D(_02947_),
    .Q(\mem_rdata_q[16] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _43104_ (.D(_02948_),
    .Q(\mem_rdata_q[17] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _43105_ (.D(_02949_),
    .Q(\mem_rdata_q[18] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _43106_ (.D(_02950_),
    .Q(\mem_rdata_q[19] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _43107_ (.D(_02951_),
    .Q(\mem_rdata_q[20] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _43108_ (.D(_02952_),
    .Q(\mem_rdata_q[21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _43109_ (.D(_02953_),
    .Q(\mem_rdata_q[22] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _43110_ (.D(_02954_),
    .Q(\mem_rdata_q[23] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_2 _43111_ (.D(_02955_),
    .Q(\mem_rdata_q[24] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43112_ (.D(_02956_),
    .Q(\mem_rdata_q[25] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_2 _43113_ (.D(_02957_),
    .Q(\mem_rdata_q[26] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_2 _43114_ (.D(_02958_),
    .Q(\mem_rdata_q[27] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _43115_ (.D(_02959_),
    .Q(\mem_rdata_q[28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43116_ (.D(_02960_),
    .Q(\mem_rdata_q[29] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _43117_ (.D(_02961_),
    .Q(\mem_rdata_q[30] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43118_ (.D(_02962_),
    .Q(\mem_rdata_q[31] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 _43119_ (.D(_02963_),
    .Q(\cpuregs[2][0] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43120_ (.D(_02964_),
    .Q(\cpuregs[2][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _43121_ (.D(_02965_),
    .Q(\cpuregs[2][2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43122_ (.D(_02966_),
    .Q(\cpuregs[2][3] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43123_ (.D(_02967_),
    .Q(\cpuregs[2][4] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43124_ (.D(_02968_),
    .Q(\cpuregs[2][5] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43125_ (.D(_02969_),
    .Q(\cpuregs[2][6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43126_ (.D(_02970_),
    .Q(\cpuregs[2][7] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43127_ (.D(_02971_),
    .Q(\cpuregs[2][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43128_ (.D(_02972_),
    .Q(\cpuregs[2][9] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43129_ (.D(_02973_),
    .Q(\cpuregs[2][10] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43130_ (.D(_02974_),
    .Q(\cpuregs[2][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43131_ (.D(_02975_),
    .Q(\cpuregs[2][12] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43132_ (.D(_02976_),
    .Q(\cpuregs[2][13] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _43133_ (.D(_02977_),
    .Q(\cpuregs[2][14] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43134_ (.D(_02978_),
    .Q(\cpuregs[2][15] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43135_ (.D(_02979_),
    .Q(\cpuregs[2][16] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43136_ (.D(_02980_),
    .Q(\cpuregs[2][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43137_ (.D(_02981_),
    .Q(\cpuregs[2][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43138_ (.D(_02982_),
    .Q(\cpuregs[2][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43139_ (.D(_02983_),
    .Q(\cpuregs[2][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43140_ (.D(_02984_),
    .Q(\cpuregs[2][21] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43141_ (.D(_02985_),
    .Q(\cpuregs[2][22] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43142_ (.D(_02986_),
    .Q(\cpuregs[2][23] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43143_ (.D(_02987_),
    .Q(\cpuregs[2][24] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43144_ (.D(_02988_),
    .Q(\cpuregs[2][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43145_ (.D(_02989_),
    .Q(\cpuregs[2][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43146_ (.D(_02990_),
    .Q(\cpuregs[2][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43147_ (.D(_02991_),
    .Q(\cpuregs[2][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43148_ (.D(_02992_),
    .Q(\cpuregs[2][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43149_ (.D(_02993_),
    .Q(\cpuregs[2][30] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43150_ (.D(_02994_),
    .Q(\cpuregs[2][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43151_ (.D(_02995_),
    .Q(\cpuregs[5][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43152_ (.D(_02996_),
    .Q(\cpuregs[5][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43153_ (.D(_02997_),
    .Q(\cpuregs[5][2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43154_ (.D(_02998_),
    .Q(\cpuregs[5][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43155_ (.D(_02999_),
    .Q(\cpuregs[5][4] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43156_ (.D(_03000_),
    .Q(\cpuregs[5][5] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43157_ (.D(_03001_),
    .Q(\cpuregs[5][6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43158_ (.D(_03002_),
    .Q(\cpuregs[5][7] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43159_ (.D(_03003_),
    .Q(\cpuregs[5][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43160_ (.D(_03004_),
    .Q(\cpuregs[5][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43161_ (.D(_03005_),
    .Q(\cpuregs[5][10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43162_ (.D(_03006_),
    .Q(\cpuregs[5][11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43163_ (.D(_03007_),
    .Q(\cpuregs[5][12] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43164_ (.D(_03008_),
    .Q(\cpuregs[5][13] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _43165_ (.D(_03009_),
    .Q(\cpuregs[5][14] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43166_ (.D(_03010_),
    .Q(\cpuregs[5][15] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43167_ (.D(_03011_),
    .Q(\cpuregs[5][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43168_ (.D(_03012_),
    .Q(\cpuregs[5][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43169_ (.D(_03013_),
    .Q(\cpuregs[5][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43170_ (.D(_03014_),
    .Q(\cpuregs[5][19] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43171_ (.D(_03015_),
    .Q(\cpuregs[5][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43172_ (.D(_03016_),
    .Q(\cpuregs[5][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43173_ (.D(_03017_),
    .Q(\cpuregs[5][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43174_ (.D(_03018_),
    .Q(\cpuregs[5][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43175_ (.D(_03019_),
    .Q(\cpuregs[5][24] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _43176_ (.D(_03020_),
    .Q(\cpuregs[5][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43177_ (.D(_03021_),
    .Q(\cpuregs[5][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43178_ (.D(_03022_),
    .Q(\cpuregs[5][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43179_ (.D(_03023_),
    .Q(\cpuregs[5][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43180_ (.D(_03024_),
    .Q(\cpuregs[5][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43181_ (.D(_03025_),
    .Q(\cpuregs[5][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43182_ (.D(_03026_),
    .Q(\cpuregs[5][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _43183_ (.D(_03027_),
    .Q(\pcpi_mul.rs1[0] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_4 _43184_ (.D(_03028_),
    .Q(\pcpi_mul.rs1[1] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_2 _43185_ (.D(_03029_),
    .Q(\pcpi_mul.rs1[2] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_4 _43186_ (.D(_03030_),
    .Q(\pcpi_mul.rs1[3] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_2 _43187_ (.D(_03031_),
    .Q(\pcpi_mul.rs1[4] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_2 _43188_ (.D(_03032_),
    .Q(\pcpi_mul.rs1[5] ),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _43189_ (.D(_03033_),
    .Q(\pcpi_mul.rs1[6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 _43190_ (.D(_03034_),
    .Q(\pcpi_mul.rs1[7] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _43191_ (.D(_03035_),
    .Q(\pcpi_mul.rs1[8] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _43192_ (.D(_03036_),
    .Q(\pcpi_mul.rs1[9] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 _43193_ (.D(_03037_),
    .Q(\pcpi_mul.rs1[10] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_1 _43194_ (.D(_03038_),
    .Q(\pcpi_mul.rs1[11] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _43195_ (.D(_03039_),
    .Q(\pcpi_mul.rs1[12] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _43196_ (.D(_03040_),
    .Q(\pcpi_mul.rs1[13] ),
    .CLK(clknet_5_26_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43197_ (.D(_03041_),
    .Q(\pcpi_mul.rs1[14] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_1 _43198_ (.D(_03042_),
    .Q(\pcpi_mul.rs1[15] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _43199_ (.D(_03043_),
    .Q(\pcpi_mul.rs1[16] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _43200_ (.D(_03044_),
    .Q(\pcpi_mul.rs1[17] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_1 _43201_ (.D(_03045_),
    .Q(\pcpi_mul.rs1[18] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 _43202_ (.D(_03046_),
    .Q(\pcpi_mul.rs1[19] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_2 _43203_ (.D(_03047_),
    .Q(\pcpi_mul.rs1[20] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_4 _43204_ (.D(_03048_),
    .Q(\pcpi_mul.rs1[21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 _43205_ (.D(_03049_),
    .Q(\pcpi_mul.rs1[22] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_2 _43206_ (.D(_03050_),
    .Q(\pcpi_mul.rs1[23] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 _43207_ (.D(_03051_),
    .Q(\pcpi_mul.rs1[24] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 _43208_ (.D(_03052_),
    .Q(\pcpi_mul.rs1[25] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_4 _43209_ (.D(_03053_),
    .Q(\pcpi_mul.rs1[26] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _43210_ (.D(_03054_),
    .Q(\pcpi_mul.rs1[27] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _43211_ (.D(_03055_),
    .Q(\pcpi_mul.rs1[28] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _43212_ (.D(_03056_),
    .Q(\pcpi_mul.rs1[29] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_4 _43213_ (.D(_03057_),
    .Q(\pcpi_mul.rs1[30] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_4 _43214_ (.D(_03058_),
    .Q(\pcpi_mul.rs1[31] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 _43215_ (.D(_03059_),
    .Q(net156),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_4 _43216_ (.D(_03060_),
    .Q(net159),
    .CLK(clknet_5_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43217_ (.D(_03061_),
    .Q(net160),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_1 _43218_ (.D(_03062_),
    .Q(net161),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_4 _43219_ (.D(_03063_),
    .Q(net162),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_4 _43220_ (.D(_03064_),
    .Q(net163),
    .CLK(clknet_opt_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43221_ (.D(_03065_),
    .Q(net164),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _43222_ (.D(_03066_),
    .Q(net165),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 _43223_ (.D(_03067_),
    .Q(net135),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 _43224_ (.D(_03068_),
    .Q(net136),
    .CLK(clknet_opt_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _43225_ (.D(_03069_),
    .Q(net137),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_1 _43226_ (.D(_03070_),
    .Q(net138),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _43227_ (.D(_03071_),
    .Q(net139),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43228_ (.D(_03072_),
    .Q(net140),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43229_ (.D(_03073_),
    .Q(net141),
    .CLK(clknet_5_30_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43230_ (.D(_03074_),
    .Q(net142),
    .CLK(clknet_opt_7_clk));
 sky130_fd_sc_hd__dfxtp_4 _43231_ (.D(_03075_),
    .Q(net143),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _43232_ (.D(_03076_),
    .Q(net144),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_4 _43233_ (.D(_03077_),
    .Q(net146),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _43234_ (.D(_03078_),
    .Q(net147),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 _43235_ (.D(_03079_),
    .Q(net148),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _43236_ (.D(_03080_),
    .Q(net149),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_4 _43237_ (.D(_03081_),
    .Q(net150),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_4 _43238_ (.D(_03082_),
    .Q(net151),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_4 _43239_ (.D(_03083_),
    .Q(net152),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_4 _43240_ (.D(_03084_),
    .Q(net153),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _43241_ (.D(_03085_),
    .Q(net154),
    .CLK(clknet_opt_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43242_ (.D(_03086_),
    .Q(net155),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_1 _43243_ (.D(_03087_),
    .Q(net157),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _43244_ (.D(_03088_),
    .Q(net158),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_4 _43245_ (.D(_03089_),
    .Q(net306),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_4 _43246_ (.D(_03090_),
    .Q(net317),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43247_ (.D(_03091_),
    .Q(net328),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_4 _43248_ (.D(_03092_),
    .Q(net331),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_4 _43249_ (.D(_03093_),
    .Q(net332),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_4 _43250_ (.D(_03094_),
    .Q(net333),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_4 _43251_ (.D(_03095_),
    .Q(net334),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_4 _43252_ (.D(_03096_),
    .Q(net335),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_4 _43253_ (.D(_03097_),
    .Q(net336),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _43254_ (.D(_03098_),
    .Q(net337),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _43255_ (.D(_03099_),
    .Q(net307),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _43256_ (.D(_03100_),
    .Q(net308),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_4 _43257_ (.D(_03101_),
    .Q(net309),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_4 _43258_ (.D(_03102_),
    .Q(net310),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_4 _43259_ (.D(_03103_),
    .Q(net311),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_4 _43260_ (.D(_03104_),
    .Q(net312),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_4 _43261_ (.D(_03105_),
    .Q(net313),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_4 _43262_ (.D(_03106_),
    .Q(net314),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_4 _43263_ (.D(_03107_),
    .Q(net315),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_4 _43264_ (.D(_03108_),
    .Q(net316),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_4 _43265_ (.D(_03109_),
    .Q(net318),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_4 _43266_ (.D(_03110_),
    .Q(net319),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_4 _43267_ (.D(_03111_),
    .Q(net320),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_4 _43268_ (.D(_03112_),
    .Q(net321),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_4 _43269_ (.D(_03113_),
    .Q(net322),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_4 _43270_ (.D(_03114_),
    .Q(net323),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43271_ (.D(_03115_),
    .Q(net324),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_4 _43272_ (.D(_03116_),
    .Q(net325),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_4 _43273_ (.D(_03117_),
    .Q(net326),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_4 _43274_ (.D(_03118_),
    .Q(net327),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_4 _43275_ (.D(_03119_),
    .Q(net329),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_4 _43276_ (.D(_03120_),
    .Q(net330),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_4 _43277_ (.D(_03121_),
    .Q(net274),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_4 _43278_ (.D(_03122_),
    .Q(net285),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _43279_ (.D(_03123_),
    .Q(net296),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _43280_ (.D(_03124_),
    .Q(net299),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_4 _43281_ (.D(_03125_),
    .Q(net300),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_4 _43282_ (.D(_03126_),
    .Q(net301),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 _43283_ (.D(_03127_),
    .Q(net302),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_4 _43284_ (.D(_03128_),
    .Q(net303),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_4 _43285_ (.D(_03129_),
    .Q(net304),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_4 _43286_ (.D(_03130_),
    .Q(net305),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _43287_ (.D(_03131_),
    .Q(net275),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _43288_ (.D(_03132_),
    .Q(net276),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_4 _43289_ (.D(_03133_),
    .Q(net277),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_4 _43290_ (.D(_03134_),
    .Q(net278),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 _43291_ (.D(_03135_),
    .Q(net279),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 _43292_ (.D(_03136_),
    .Q(net280),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _43293_ (.D(_03137_),
    .Q(net281),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _43294_ (.D(_03138_),
    .Q(net282),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _43295_ (.D(_03139_),
    .Q(net283),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _43296_ (.D(_03140_),
    .Q(net284),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_4 _43297_ (.D(_03141_),
    .Q(net286),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _43298_ (.D(_03142_),
    .Q(net287),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _43299_ (.D(_03143_),
    .Q(net288),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _43300_ (.D(_03144_),
    .Q(net289),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _43301_ (.D(_03145_),
    .Q(net290),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_4 _43302_ (.D(_03146_),
    .Q(net291),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_2 _43303_ (.D(_03147_),
    .Q(net292),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_4 _43304_ (.D(_03148_),
    .Q(net293),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_4 _43305_ (.D(_03149_),
    .Q(net294),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_4 _43306_ (.D(_03150_),
    .Q(net295),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_2 _43307_ (.D(_03151_),
    .Q(net297),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_4 _43308_ (.D(_03152_),
    .Q(net298),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_4 _43309_ (.D(_03153_),
    .Q(instr_lui),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_2 _43310_ (.D(_03154_),
    .Q(instr_auipc),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_4 _43311_ (.D(_03155_),
    .Q(instr_jal),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 _43312_ (.D(_03156_),
    .Q(instr_jalr),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43313_ (.D(_03157_),
    .Q(instr_lb),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43314_ (.D(_03158_),
    .Q(instr_lh),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43315_ (.D(_03159_),
    .Q(instr_lw),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43316_ (.D(_03160_),
    .Q(instr_lbu),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43317_ (.D(_03161_),
    .Q(instr_lhu),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43318_ (.D(_03162_),
    .Q(instr_sb),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43319_ (.D(_03163_),
    .Q(instr_sh),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43320_ (.D(_03164_),
    .Q(instr_sw),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_2 _43321_ (.D(_03165_),
    .Q(instr_slli),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43322_ (.D(_03166_),
    .Q(instr_srli),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _43323_ (.D(_03167_),
    .Q(instr_srai),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _43324_ (.D(_03168_),
    .Q(instr_rdcycle),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_2 _43325_ (.D(_03169_),
    .Q(instr_rdcycleh),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43326_ (.D(_03170_),
    .Q(instr_rdinstr),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43327_ (.D(_03171_),
    .Q(instr_rdinstrh),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43328_ (.D(_03172_),
    .Q(instr_ecall_ebreak),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43329_ (.D(_03173_),
    .Q(instr_getq),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_2 _43330_ (.D(_03174_),
    .Q(instr_setq),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43331_ (.D(_03175_),
    .Q(instr_retirq),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43332_ (.D(_03176_),
    .Q(instr_maskirq),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_2 _43333_ (.D(_03177_),
    .Q(instr_waitirq),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_4 _43334_ (.D(_03178_),
    .Q(instr_timer),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43335_ (.D(_03179_),
    .Q(\decoded_rd[0] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _43336_ (.D(_03180_),
    .Q(\decoded_rd[1] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_4 _43337_ (.D(_03181_),
    .Q(\decoded_rd[2] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_4 _43338_ (.D(_03182_),
    .Q(\decoded_rd[3] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 _43339_ (.D(_03183_),
    .Q(\decoded_rd[4] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _43340_ (.D(_03184_),
    .Q(\decoded_imm[0] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_2 _43341_ (.D(_03185_),
    .Q(\decoded_imm_uj[1] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _43342_ (.D(_03186_),
    .Q(\decoded_imm_uj[2] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _43343_ (.D(_03187_),
    .Q(\decoded_imm_uj[3] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _43344_ (.D(_03188_),
    .Q(\decoded_imm_uj[4] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43345_ (.D(_03189_),
    .Q(\decoded_imm_uj[5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43346_ (.D(_03190_),
    .Q(\decoded_imm_uj[6] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43347_ (.D(_03191_),
    .Q(\decoded_imm_uj[7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _43348_ (.D(_03192_),
    .Q(\decoded_imm_uj[8] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43349_ (.D(_03193_),
    .Q(\decoded_imm_uj[9] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _43350_ (.D(_03194_),
    .Q(\decoded_imm_uj[10] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_4 _43351_ (.D(_03195_),
    .Q(\decoded_imm_uj[11] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _43352_ (.D(_03196_),
    .Q(\decoded_imm_uj[12] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _43353_ (.D(_03197_),
    .Q(\decoded_imm_uj[13] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _43354_ (.D(_03198_),
    .Q(\decoded_imm_uj[14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_4 _43355_ (.D(_03199_),
    .Q(\decoded_imm_uj[15] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_4 _43356_ (.D(_03200_),
    .Q(\decoded_imm_uj[16] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_4 _43357_ (.D(_03201_),
    .Q(\decoded_imm_uj[17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_4 _43358_ (.D(_03202_),
    .Q(\decoded_imm_uj[18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_4 _43359_ (.D(_03203_),
    .Q(\decoded_imm_uj[19] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_2 _43360_ (.D(_03204_),
    .Q(\decoded_imm_uj[20] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43361_ (.D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_4 _43362_ (.D(_03206_),
    .Q(is_slli_srli_srai),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43363_ (.D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43364_ (.D(_03208_),
    .Q(is_sb_sh_sw),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43365_ (.D(_03209_),
    .Q(\cpuregs[13][0] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43366_ (.D(_03210_),
    .Q(\cpuregs[13][1] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _43367_ (.D(_03211_),
    .Q(\cpuregs[13][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43368_ (.D(_03212_),
    .Q(\cpuregs[13][3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43369_ (.D(_03213_),
    .Q(\cpuregs[13][4] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43370_ (.D(_03214_),
    .Q(\cpuregs[13][5] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43371_ (.D(_03215_),
    .Q(\cpuregs[13][6] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43372_ (.D(_03216_),
    .Q(\cpuregs[13][7] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43373_ (.D(_03217_),
    .Q(\cpuregs[13][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43374_ (.D(_03218_),
    .Q(\cpuregs[13][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43375_ (.D(_03219_),
    .Q(\cpuregs[13][10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43376_ (.D(_03220_),
    .Q(\cpuregs[13][11] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _43377_ (.D(_03221_),
    .Q(\cpuregs[13][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43378_ (.D(_03222_),
    .Q(\cpuregs[13][13] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 _43379_ (.D(_03223_),
    .Q(\cpuregs[13][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43380_ (.D(_03224_),
    .Q(\cpuregs[13][15] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43381_ (.D(_03225_),
    .Q(\cpuregs[13][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43382_ (.D(_03226_),
    .Q(\cpuregs[13][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43383_ (.D(_03227_),
    .Q(\cpuregs[13][18] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43384_ (.D(_03228_),
    .Q(\cpuregs[13][19] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43385_ (.D(_03229_),
    .Q(\cpuregs[13][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43386_ (.D(_03230_),
    .Q(\cpuregs[13][21] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43387_ (.D(_03231_),
    .Q(\cpuregs[13][22] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _43388_ (.D(_03232_),
    .Q(\cpuregs[13][23] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _43389_ (.D(_03233_),
    .Q(\cpuregs[13][24] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _43390_ (.D(_03234_),
    .Q(\cpuregs[13][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43391_ (.D(_03235_),
    .Q(\cpuregs[13][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43392_ (.D(_03236_),
    .Q(\cpuregs[13][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43393_ (.D(_03237_),
    .Q(\cpuregs[13][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43394_ (.D(_03238_),
    .Q(\cpuregs[13][29] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43395_ (.D(_03239_),
    .Q(\cpuregs[13][30] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43396_ (.D(_03240_),
    .Q(\cpuregs[13][31] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43397_ (.D(_03241_),
    .Q(is_alu_reg_imm),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _43398_ (.D(_03242_),
    .Q(is_alu_reg_reg),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_4 _43399_ (.D(_03243_),
    .Q(net270),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_4 _43400_ (.D(_03244_),
    .Q(net271),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_4 _43401_ (.D(_03245_),
    .Q(net272),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_4 _43402_ (.D(_03246_),
    .Q(net273),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _43403_ (.D(_03247_),
    .Q(\pcpi_mul.rs2[0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_1 _43404_ (.D(_03248_),
    .Q(\pcpi_mul.rs2[1] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _43405_ (.D(_03249_),
    .Q(\pcpi_mul.rs2[2] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _43406_ (.D(_03250_),
    .Q(\pcpi_mul.rs2[3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43407_ (.D(_03251_),
    .Q(\pcpi_mul.rs2[4] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _43408_ (.D(_03252_),
    .Q(\pcpi_mul.rs2[5] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_2 _43409_ (.D(_03253_),
    .Q(\pcpi_mul.rs2[6] ),
    .CLK(clknet_5_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43410_ (.D(_03254_),
    .Q(\pcpi_mul.rs2[7] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _43411_ (.D(_03255_),
    .Q(\pcpi_mul.rs2[8] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_1 _43412_ (.D(_03256_),
    .Q(\pcpi_mul.rs2[9] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 _43413_ (.D(_03257_),
    .Q(\pcpi_mul.rs2[10] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 _43414_ (.D(_03258_),
    .Q(\pcpi_mul.rs2[11] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _43415_ (.D(_03259_),
    .Q(\pcpi_mul.rs2[12] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_4 _43416_ (.D(_03260_),
    .Q(\pcpi_mul.rs2[13] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _43417_ (.D(_03261_),
    .Q(\pcpi_mul.rs2[14] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 _43418_ (.D(_03262_),
    .Q(\pcpi_mul.rs2[15] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_1 _43419_ (.D(_03263_),
    .Q(\pcpi_mul.rs2[16] ),
    .CLK(clknet_5_26_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _43420_ (.D(_03264_),
    .Q(\pcpi_mul.rs2[17] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43421_ (.D(_03265_),
    .Q(\pcpi_mul.rs2[18] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _43422_ (.D(_03266_),
    .Q(\pcpi_mul.rs2[19] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_4 _43423_ (.D(_03267_),
    .Q(\pcpi_mul.rs2[20] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_4 _43424_ (.D(_03268_),
    .Q(\pcpi_mul.rs2[21] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_4 _43425_ (.D(_03269_),
    .Q(\pcpi_mul.rs2[22] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _43426_ (.D(_03270_),
    .Q(\pcpi_mul.rs2[23] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_4 _43427_ (.D(_03271_),
    .Q(\pcpi_mul.rs2[24] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_2 _43428_ (.D(_03272_),
    .Q(\pcpi_mul.rs2[25] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_2 _43429_ (.D(_03273_),
    .Q(\pcpi_mul.rs2[26] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_4 _43430_ (.D(_03274_),
    .Q(\pcpi_mul.rs2[27] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_4 _43431_ (.D(_03275_),
    .Q(\pcpi_mul.rs2[28] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_4 _43432_ (.D(_03276_),
    .Q(\pcpi_mul.rs2[29] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_2 _43433_ (.D(_03277_),
    .Q(\pcpi_mul.rs2[30] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _43434_ (.D(_03278_),
    .Q(\pcpi_mul.rs2[31] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 _43435_ (.D(_03279_),
    .Q(\cpuregs[17][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43436_ (.D(_03280_),
    .Q(\cpuregs[17][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43437_ (.D(_03281_),
    .Q(\cpuregs[17][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43438_ (.D(_03282_),
    .Q(\cpuregs[17][3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43439_ (.D(_03283_),
    .Q(\cpuregs[17][4] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43440_ (.D(_03284_),
    .Q(\cpuregs[17][5] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43441_ (.D(_03285_),
    .Q(\cpuregs[17][6] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43442_ (.D(_03286_),
    .Q(\cpuregs[17][7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43443_ (.D(_03287_),
    .Q(\cpuregs[17][8] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43444_ (.D(_03288_),
    .Q(\cpuregs[17][9] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43445_ (.D(_03289_),
    .Q(\cpuregs[17][10] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43446_ (.D(_03290_),
    .Q(\cpuregs[17][11] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43447_ (.D(_03291_),
    .Q(\cpuregs[17][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43448_ (.D(_03292_),
    .Q(\cpuregs[17][13] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43449_ (.D(_03293_),
    .Q(\cpuregs[17][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43450_ (.D(_03294_),
    .Q(\cpuregs[17][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43451_ (.D(_03295_),
    .Q(\cpuregs[17][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43452_ (.D(_03296_),
    .Q(\cpuregs[17][17] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43453_ (.D(_03297_),
    .Q(\cpuregs[17][18] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43454_ (.D(_03298_),
    .Q(\cpuregs[17][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43455_ (.D(_03299_),
    .Q(\cpuregs[17][20] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _43456_ (.D(_03300_),
    .Q(\cpuregs[17][21] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_1 _43457_ (.D(_03301_),
    .Q(\cpuregs[17][22] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43458_ (.D(_03302_),
    .Q(\cpuregs[17][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43459_ (.D(_03303_),
    .Q(\cpuregs[17][24] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _43460_ (.D(_03304_),
    .Q(\cpuregs[17][25] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43461_ (.D(_03305_),
    .Q(\cpuregs[17][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43462_ (.D(_03306_),
    .Q(\cpuregs[17][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43463_ (.D(_03307_),
    .Q(\cpuregs[17][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43464_ (.D(_03308_),
    .Q(\cpuregs[17][29] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43465_ (.D(_03309_),
    .Q(\cpuregs[17][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43466_ (.D(_03310_),
    .Q(\cpuregs[17][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43467_ (.D(_03311_),
    .Q(\cpuregs[16][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43468_ (.D(_03312_),
    .Q(\cpuregs[16][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43469_ (.D(_03313_),
    .Q(\cpuregs[16][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43470_ (.D(_03314_),
    .Q(\cpuregs[16][3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43471_ (.D(_03315_),
    .Q(\cpuregs[16][4] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43472_ (.D(_03316_),
    .Q(\cpuregs[16][5] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43473_ (.D(_03317_),
    .Q(\cpuregs[16][6] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43474_ (.D(_03318_),
    .Q(\cpuregs[16][7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43475_ (.D(_03319_),
    .Q(\cpuregs[16][8] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 _43476_ (.D(_03320_),
    .Q(\cpuregs[16][9] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43477_ (.D(_03321_),
    .Q(\cpuregs[16][10] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43478_ (.D(_03322_),
    .Q(\cpuregs[16][11] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43479_ (.D(_03323_),
    .Q(\cpuregs[16][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43480_ (.D(_03324_),
    .Q(\cpuregs[16][13] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43481_ (.D(_03325_),
    .Q(\cpuregs[16][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43482_ (.D(_03326_),
    .Q(\cpuregs[16][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43483_ (.D(_03327_),
    .Q(\cpuregs[16][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43484_ (.D(_03328_),
    .Q(\cpuregs[16][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43485_ (.D(_03329_),
    .Q(\cpuregs[16][18] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43486_ (.D(_03330_),
    .Q(\cpuregs[16][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43487_ (.D(_03331_),
    .Q(\cpuregs[16][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43488_ (.D(_03332_),
    .Q(\cpuregs[16][21] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43489_ (.D(_03333_),
    .Q(\cpuregs[16][22] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _43490_ (.D(_03334_),
    .Q(\cpuregs[16][23] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _43491_ (.D(_03335_),
    .Q(\cpuregs[16][24] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _43492_ (.D(_03336_),
    .Q(\cpuregs[16][25] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43493_ (.D(_03337_),
    .Q(\cpuregs[16][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43494_ (.D(_03338_),
    .Q(\cpuregs[16][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43495_ (.D(_03339_),
    .Q(\cpuregs[16][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43496_ (.D(_03340_),
    .Q(\cpuregs[16][29] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43497_ (.D(_03341_),
    .Q(\cpuregs[16][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43498_ (.D(_03342_),
    .Q(\cpuregs[16][31] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _43499_ (.D(_03343_),
    .Q(\cpuregs[12][0] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43500_ (.D(_03344_),
    .Q(\cpuregs[12][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _43501_ (.D(_03345_),
    .Q(\cpuregs[12][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43502_ (.D(_03346_),
    .Q(\cpuregs[12][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43503_ (.D(_03347_),
    .Q(\cpuregs[12][4] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43504_ (.D(_03348_),
    .Q(\cpuregs[12][5] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43505_ (.D(_03349_),
    .Q(\cpuregs[12][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43506_ (.D(_03350_),
    .Q(\cpuregs[12][7] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43507_ (.D(_03351_),
    .Q(\cpuregs[12][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43508_ (.D(_03352_),
    .Q(\cpuregs[12][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43509_ (.D(_03353_),
    .Q(\cpuregs[12][10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43510_ (.D(_03354_),
    .Q(\cpuregs[12][11] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _43511_ (.D(_03355_),
    .Q(\cpuregs[12][12] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43512_ (.D(_03356_),
    .Q(\cpuregs[12][13] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _43513_ (.D(_03357_),
    .Q(\cpuregs[12][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43514_ (.D(_03358_),
    .Q(\cpuregs[12][15] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43515_ (.D(_03359_),
    .Q(\cpuregs[12][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43516_ (.D(_03360_),
    .Q(\cpuregs[12][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43517_ (.D(_03361_),
    .Q(\cpuregs[12][18] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _43518_ (.D(_03362_),
    .Q(\cpuregs[12][19] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _43519_ (.D(_03363_),
    .Q(\cpuregs[12][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43520_ (.D(_03364_),
    .Q(\cpuregs[12][21] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43521_ (.D(_03365_),
    .Q(\cpuregs[12][22] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _43522_ (.D(_03366_),
    .Q(\cpuregs[12][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43523_ (.D(_03367_),
    .Q(\cpuregs[12][24] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _43524_ (.D(_03368_),
    .Q(\cpuregs[12][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43525_ (.D(_03369_),
    .Q(\cpuregs[12][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43526_ (.D(_03370_),
    .Q(\cpuregs[12][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43527_ (.D(_03371_),
    .Q(\cpuregs[12][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43528_ (.D(_03372_),
    .Q(\cpuregs[12][29] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43529_ (.D(_03373_),
    .Q(\cpuregs[12][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43530_ (.D(_03374_),
    .Q(\cpuregs[12][31] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43531_ (.D(_03375_),
    .Q(\cpuregs[1][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43532_ (.D(_03376_),
    .Q(\cpuregs[1][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _43533_ (.D(_03377_),
    .Q(\cpuregs[1][2] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _43534_ (.D(_03378_),
    .Q(\cpuregs[1][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43535_ (.D(_03379_),
    .Q(\cpuregs[1][4] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43536_ (.D(_03380_),
    .Q(\cpuregs[1][5] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43537_ (.D(_03381_),
    .Q(\cpuregs[1][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43538_ (.D(_03382_),
    .Q(\cpuregs[1][7] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43539_ (.D(_03383_),
    .Q(\cpuregs[1][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43540_ (.D(_03384_),
    .Q(\cpuregs[1][9] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43541_ (.D(_03385_),
    .Q(\cpuregs[1][10] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43542_ (.D(_03386_),
    .Q(\cpuregs[1][11] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43543_ (.D(_03387_),
    .Q(\cpuregs[1][12] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43544_ (.D(_03388_),
    .Q(\cpuregs[1][13] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _43545_ (.D(_03389_),
    .Q(\cpuregs[1][14] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43546_ (.D(_03390_),
    .Q(\cpuregs[1][15] ),
    .CLK(clknet_5_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43547_ (.D(_03391_),
    .Q(\cpuregs[1][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43548_ (.D(_03392_),
    .Q(\cpuregs[1][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43549_ (.D(_03393_),
    .Q(\cpuregs[1][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43550_ (.D(_03394_),
    .Q(\cpuregs[1][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43551_ (.D(_03395_),
    .Q(\cpuregs[1][20] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43552_ (.D(_03396_),
    .Q(\cpuregs[1][21] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43553_ (.D(_03397_),
    .Q(\cpuregs[1][22] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43554_ (.D(_03398_),
    .Q(\cpuregs[1][23] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _43555_ (.D(_03399_),
    .Q(\cpuregs[1][24] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _43556_ (.D(_03400_),
    .Q(\cpuregs[1][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43557_ (.D(_03401_),
    .Q(\cpuregs[1][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43558_ (.D(_03402_),
    .Q(\cpuregs[1][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43559_ (.D(_03403_),
    .Q(\cpuregs[1][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43560_ (.D(_03404_),
    .Q(\cpuregs[1][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43561_ (.D(_03405_),
    .Q(\cpuregs[1][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43562_ (.D(_03406_),
    .Q(\cpuregs[1][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43563_ (.D(_03407_),
    .Q(\cpuregs[3][0] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43564_ (.D(_03408_),
    .Q(\cpuregs[3][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _43565_ (.D(_03409_),
    .Q(\cpuregs[3][2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43566_ (.D(_03410_),
    .Q(\cpuregs[3][3] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43567_ (.D(_03411_),
    .Q(\cpuregs[3][4] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43568_ (.D(_03412_),
    .Q(\cpuregs[3][5] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43569_ (.D(_03413_),
    .Q(\cpuregs[3][6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43570_ (.D(_03414_),
    .Q(\cpuregs[3][7] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43571_ (.D(_03415_),
    .Q(\cpuregs[3][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43572_ (.D(_03416_),
    .Q(\cpuregs[3][9] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43573_ (.D(_03417_),
    .Q(\cpuregs[3][10] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43574_ (.D(_03418_),
    .Q(\cpuregs[3][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43575_ (.D(_03419_),
    .Q(\cpuregs[3][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43576_ (.D(_03420_),
    .Q(\cpuregs[3][13] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _43577_ (.D(_03421_),
    .Q(\cpuregs[3][14] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43578_ (.D(_03422_),
    .Q(\cpuregs[3][15] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43579_ (.D(_03423_),
    .Q(\cpuregs[3][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43580_ (.D(_03424_),
    .Q(\cpuregs[3][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43581_ (.D(_03425_),
    .Q(\cpuregs[3][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43582_ (.D(_03426_),
    .Q(\cpuregs[3][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43583_ (.D(_03427_),
    .Q(\cpuregs[3][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43584_ (.D(_03428_),
    .Q(\cpuregs[3][21] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43585_ (.D(_03429_),
    .Q(\cpuregs[3][22] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_1 _43586_ (.D(_03430_),
    .Q(\cpuregs[3][23] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43587_ (.D(_03431_),
    .Q(\cpuregs[3][24] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _43588_ (.D(_03432_),
    .Q(\cpuregs[3][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43589_ (.D(_03433_),
    .Q(\cpuregs[3][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43590_ (.D(_03434_),
    .Q(\cpuregs[3][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43591_ (.D(_03435_),
    .Q(\cpuregs[3][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43592_ (.D(_03436_),
    .Q(\cpuregs[3][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43593_ (.D(_03437_),
    .Q(\cpuregs[3][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43594_ (.D(_03438_),
    .Q(\cpuregs[3][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43595_ (.D(_03439_),
    .Q(\cpuregs[11][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43596_ (.D(_03440_),
    .Q(\cpuregs[11][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43597_ (.D(_03441_),
    .Q(\cpuregs[11][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43598_ (.D(_03442_),
    .Q(\cpuregs[11][3] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43599_ (.D(_03443_),
    .Q(\cpuregs[11][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43600_ (.D(_03444_),
    .Q(\cpuregs[11][5] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43601_ (.D(_03445_),
    .Q(\cpuregs[11][6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43602_ (.D(_03446_),
    .Q(\cpuregs[11][7] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43603_ (.D(_03447_),
    .Q(\cpuregs[11][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43604_ (.D(_03448_),
    .Q(\cpuregs[11][9] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43605_ (.D(_03449_),
    .Q(\cpuregs[11][10] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43606_ (.D(_03450_),
    .Q(\cpuregs[11][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43607_ (.D(_03451_),
    .Q(\cpuregs[11][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43608_ (.D(_03452_),
    .Q(\cpuregs[11][13] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43609_ (.D(_03453_),
    .Q(\cpuregs[11][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43610_ (.D(_03454_),
    .Q(\cpuregs[11][15] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43611_ (.D(_03455_),
    .Q(\cpuregs[11][16] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43612_ (.D(_03456_),
    .Q(\cpuregs[11][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43613_ (.D(_03457_),
    .Q(\cpuregs[11][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43614_ (.D(_03458_),
    .Q(\cpuregs[11][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43615_ (.D(_03459_),
    .Q(\cpuregs[11][20] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43616_ (.D(_03460_),
    .Q(\cpuregs[11][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43617_ (.D(_03461_),
    .Q(\cpuregs[11][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43618_ (.D(_03462_),
    .Q(\cpuregs[11][23] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _43619_ (.D(_03463_),
    .Q(\cpuregs[11][24] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _43620_ (.D(_03464_),
    .Q(\cpuregs[11][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43621_ (.D(_03465_),
    .Q(\cpuregs[11][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43622_ (.D(_03466_),
    .Q(\cpuregs[11][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43623_ (.D(_03467_),
    .Q(\cpuregs[11][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43624_ (.D(_03468_),
    .Q(\cpuregs[11][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43625_ (.D(_03469_),
    .Q(\cpuregs[11][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43626_ (.D(_03470_),
    .Q(\cpuregs[11][31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43627_ (.D(_03471_),
    .Q(\cpuregs[15][0] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43628_ (.D(_03472_),
    .Q(\cpuregs[15][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _43629_ (.D(_03473_),
    .Q(\cpuregs[15][2] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43630_ (.D(_03474_),
    .Q(\cpuregs[15][3] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43631_ (.D(_03475_),
    .Q(\cpuregs[15][4] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43632_ (.D(_03476_),
    .Q(\cpuregs[15][5] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43633_ (.D(_03477_),
    .Q(\cpuregs[15][6] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43634_ (.D(_03478_),
    .Q(\cpuregs[15][7] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43635_ (.D(_03479_),
    .Q(\cpuregs[15][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43636_ (.D(_03480_),
    .Q(\cpuregs[15][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43637_ (.D(_03481_),
    .Q(\cpuregs[15][10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43638_ (.D(_03482_),
    .Q(\cpuregs[15][11] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43639_ (.D(_03483_),
    .Q(\cpuregs[15][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43640_ (.D(_03484_),
    .Q(\cpuregs[15][13] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _43641_ (.D(_03485_),
    .Q(\cpuregs[15][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43642_ (.D(_03486_),
    .Q(\cpuregs[15][15] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43643_ (.D(_03487_),
    .Q(\cpuregs[15][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43644_ (.D(_03488_),
    .Q(\cpuregs[15][17] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43645_ (.D(_03489_),
    .Q(\cpuregs[15][18] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43646_ (.D(_03490_),
    .Q(\cpuregs[15][19] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _43647_ (.D(_03491_),
    .Q(\cpuregs[15][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43648_ (.D(_03492_),
    .Q(\cpuregs[15][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43649_ (.D(_03493_),
    .Q(\cpuregs[15][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43650_ (.D(_03494_),
    .Q(\cpuregs[15][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43651_ (.D(_03495_),
    .Q(\cpuregs[15][24] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _43652_ (.D(_03496_),
    .Q(\cpuregs[15][25] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43653_ (.D(_03497_),
    .Q(\cpuregs[15][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43654_ (.D(_03498_),
    .Q(\cpuregs[15][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43655_ (.D(_03499_),
    .Q(\cpuregs[15][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43656_ (.D(_03500_),
    .Q(\cpuregs[15][29] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43657_ (.D(_03501_),
    .Q(\cpuregs[15][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43658_ (.D(_03502_),
    .Q(\cpuregs[15][31] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_4 _43659_ (.D(_03503_),
    .Q(\latched_rd[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _43660_ (.D(_03504_),
    .Q(\cpuregs[7][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43661_ (.D(_03505_),
    .Q(\cpuregs[7][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43662_ (.D(_03506_),
    .Q(\cpuregs[7][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43663_ (.D(_03507_),
    .Q(\cpuregs[7][3] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43664_ (.D(_03508_),
    .Q(\cpuregs[7][4] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43665_ (.D(_03509_),
    .Q(\cpuregs[7][5] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43666_ (.D(_03510_),
    .Q(\cpuregs[7][6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43667_ (.D(_03511_),
    .Q(\cpuregs[7][7] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43668_ (.D(_03512_),
    .Q(\cpuregs[7][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43669_ (.D(_03513_),
    .Q(\cpuregs[7][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43670_ (.D(_03514_),
    .Q(\cpuregs[7][10] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43671_ (.D(_03515_),
    .Q(\cpuregs[7][11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43672_ (.D(_03516_),
    .Q(\cpuregs[7][12] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43673_ (.D(_03517_),
    .Q(\cpuregs[7][13] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43674_ (.D(_03518_),
    .Q(\cpuregs[7][14] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43675_ (.D(_03519_),
    .Q(\cpuregs[7][15] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43676_ (.D(_03520_),
    .Q(\cpuregs[7][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43677_ (.D(_03521_),
    .Q(\cpuregs[7][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43678_ (.D(_03522_),
    .Q(\cpuregs[7][18] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43679_ (.D(_03523_),
    .Q(\cpuregs[7][19] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43680_ (.D(_03524_),
    .Q(\cpuregs[7][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43681_ (.D(_03525_),
    .Q(\cpuregs[7][21] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43682_ (.D(_03526_),
    .Q(\cpuregs[7][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43683_ (.D(_03527_),
    .Q(\cpuregs[7][23] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43684_ (.D(_03528_),
    .Q(\cpuregs[7][24] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43685_ (.D(_03529_),
    .Q(\cpuregs[7][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43686_ (.D(_03530_),
    .Q(\cpuregs[7][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43687_ (.D(_03531_),
    .Q(\cpuregs[7][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43688_ (.D(_03532_),
    .Q(\cpuregs[7][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43689_ (.D(_03533_),
    .Q(\cpuregs[7][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43690_ (.D(_03534_),
    .Q(\cpuregs[7][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43691_ (.D(_03535_),
    .Q(\cpuregs[7][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_4 _43692_ (.D(_03536_),
    .Q(net238),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_4 _43693_ (.D(_03537_),
    .Q(net249),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 _43694_ (.D(_03538_),
    .Q(net260),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_4 _43695_ (.D(_03539_),
    .Q(net263),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 _43696_ (.D(_03540_),
    .Q(net264),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_4 _43697_ (.D(_03541_),
    .Q(net265),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _43698_ (.D(_03542_),
    .Q(net266),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 _43699_ (.D(_03543_),
    .Q(net267),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_1 _43700_ (.D(_03544_),
    .Q(net268),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43701_ (.D(_03545_),
    .Q(net269),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _43702_ (.D(_03546_),
    .Q(net239),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _43703_ (.D(_03547_),
    .Q(net240),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_4 _43704_ (.D(_03548_),
    .Q(net241),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 _43705_ (.D(_03549_),
    .Q(net242),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43706_ (.D(_03550_),
    .Q(net243),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 _43707_ (.D(_03551_),
    .Q(net244),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43708_ (.D(_03552_),
    .Q(net245),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43709_ (.D(_03553_),
    .Q(net246),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _43710_ (.D(_03554_),
    .Q(net247),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _43711_ (.D(_03555_),
    .Q(net248),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_4 _43712_ (.D(_03556_),
    .Q(net250),
    .CLK(clknet_5_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _43713_ (.D(_03557_),
    .Q(net251),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 _43714_ (.D(_03558_),
    .Q(net252),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 _43715_ (.D(_03559_),
    .Q(net253),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 _43716_ (.D(_03560_),
    .Q(net254),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 _43717_ (.D(_03561_),
    .Q(net255),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 _43718_ (.D(_03562_),
    .Q(net256),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_4 _43719_ (.D(_03563_),
    .Q(net257),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_4 _43720_ (.D(_03564_),
    .Q(net258),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _43721_ (.D(_03565_),
    .Q(net259),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _43722_ (.D(_03566_),
    .Q(net261),
    .CLK(clknet_5_31_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _43723_ (.D(_03567_),
    .Q(net262),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 _43724_ (.D(_03568_),
    .Q(\cpuregs[19][0] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43725_ (.D(_03569_),
    .Q(\cpuregs[19][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43726_ (.D(_03570_),
    .Q(\cpuregs[19][2] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43727_ (.D(_03571_),
    .Q(\cpuregs[19][3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43728_ (.D(_03572_),
    .Q(\cpuregs[19][4] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43729_ (.D(_03573_),
    .Q(\cpuregs[19][5] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43730_ (.D(_03574_),
    .Q(\cpuregs[19][6] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43731_ (.D(_03575_),
    .Q(\cpuregs[19][7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43732_ (.D(_03576_),
    .Q(\cpuregs[19][8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43733_ (.D(_03577_),
    .Q(\cpuregs[19][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43734_ (.D(_03578_),
    .Q(\cpuregs[19][10] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43735_ (.D(_03579_),
    .Q(\cpuregs[19][11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43736_ (.D(_03580_),
    .Q(\cpuregs[19][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43737_ (.D(_03581_),
    .Q(\cpuregs[19][13] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _43738_ (.D(_03582_),
    .Q(\cpuregs[19][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43739_ (.D(_03583_),
    .Q(\cpuregs[19][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43740_ (.D(_03584_),
    .Q(\cpuregs[19][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43741_ (.D(_03585_),
    .Q(\cpuregs[19][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43742_ (.D(_03586_),
    .Q(\cpuregs[19][18] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__dfxtp_1 _43743_ (.D(_03587_),
    .Q(\cpuregs[19][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43744_ (.D(_03588_),
    .Q(\cpuregs[19][20] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43745_ (.D(_03589_),
    .Q(\cpuregs[19][21] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43746_ (.D(_03590_),
    .Q(\cpuregs[19][22] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _43747_ (.D(_03591_),
    .Q(\cpuregs[19][23] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _43748_ (.D(_03592_),
    .Q(\cpuregs[19][24] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _43749_ (.D(_03593_),
    .Q(\cpuregs[19][25] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43750_ (.D(_03594_),
    .Q(\cpuregs[19][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43751_ (.D(_03595_),
    .Q(\cpuregs[19][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43752_ (.D(_03596_),
    .Q(\cpuregs[19][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43753_ (.D(_03597_),
    .Q(\cpuregs[19][29] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43754_ (.D(_03598_),
    .Q(\cpuregs[19][30] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43755_ (.D(_03599_),
    .Q(\cpuregs[19][31] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _43756_ (.D(_03600_),
    .Q(\cpuregs[4][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43757_ (.D(_03601_),
    .Q(\cpuregs[4][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43758_ (.D(_03602_),
    .Q(\cpuregs[4][2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _43759_ (.D(_03603_),
    .Q(\cpuregs[4][3] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43760_ (.D(_03604_),
    .Q(\cpuregs[4][4] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43761_ (.D(_03605_),
    .Q(\cpuregs[4][5] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43762_ (.D(_03606_),
    .Q(\cpuregs[4][6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43763_ (.D(_03607_),
    .Q(\cpuregs[4][7] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43764_ (.D(_03608_),
    .Q(\cpuregs[4][8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43765_ (.D(_03609_),
    .Q(\cpuregs[4][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43766_ (.D(_03610_),
    .Q(\cpuregs[4][10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43767_ (.D(_03611_),
    .Q(\cpuregs[4][11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43768_ (.D(_03612_),
    .Q(\cpuregs[4][12] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43769_ (.D(_03613_),
    .Q(\cpuregs[4][13] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43770_ (.D(_03614_),
    .Q(\cpuregs[4][14] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43771_ (.D(_03615_),
    .Q(\cpuregs[4][15] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43772_ (.D(_03616_),
    .Q(\cpuregs[4][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43773_ (.D(_03617_),
    .Q(\cpuregs[4][17] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43774_ (.D(_03618_),
    .Q(\cpuregs[4][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43775_ (.D(_03619_),
    .Q(\cpuregs[4][19] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43776_ (.D(_03620_),
    .Q(\cpuregs[4][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43777_ (.D(_03621_),
    .Q(\cpuregs[4][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43778_ (.D(_03622_),
    .Q(\cpuregs[4][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43779_ (.D(_03623_),
    .Q(\cpuregs[4][23] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43780_ (.D(_03624_),
    .Q(\cpuregs[4][24] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43781_ (.D(_03625_),
    .Q(\cpuregs[4][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43782_ (.D(_03626_),
    .Q(\cpuregs[4][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43783_ (.D(_03627_),
    .Q(\cpuregs[4][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43784_ (.D(_03628_),
    .Q(\cpuregs[4][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43785_ (.D(_03629_),
    .Q(\cpuregs[4][29] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43786_ (.D(_03630_),
    .Q(\cpuregs[4][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43787_ (.D(_03631_),
    .Q(\cpuregs[4][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_4 _43788_ (.D(_03632_),
    .Q(net200),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43789_ (.D(_03633_),
    .Q(net211),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43790_ (.D(_03634_),
    .Q(net222),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43791_ (.D(_03635_),
    .Q(net225),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43792_ (.D(_03636_),
    .Q(net226),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43793_ (.D(_03637_),
    .Q(net227),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_4 _43794_ (.D(_03638_),
    .Q(net228),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_4 _43795_ (.D(_03639_),
    .Q(net229),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_4 _43796_ (.D(_03640_),
    .Q(net368),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_4 _43797_ (.D(_03641_),
    .Q(net369),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_4 _43798_ (.D(_03642_),
    .Q(net339),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _43799_ (.D(_03643_),
    .Q(net340),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_4 _43800_ (.D(_03644_),
    .Q(net341),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_4 _43801_ (.D(_03645_),
    .Q(net342),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_4 _43802_ (.D(_03646_),
    .Q(net343),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_4 _43803_ (.D(_03647_),
    .Q(net344),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_4 _43804_ (.D(_03648_),
    .Q(net345),
    .CLK(clknet_5_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _43805_ (.D(_03649_),
    .Q(net346),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_4 _43806_ (.D(_03650_),
    .Q(net347),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43807_ (.D(_03651_),
    .Q(net348),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_4 _43808_ (.D(_03652_),
    .Q(net350),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_4 _43809_ (.D(_03653_),
    .Q(net351),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43810_ (.D(_03654_),
    .Q(net352),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43811_ (.D(_03655_),
    .Q(net353),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43812_ (.D(_03656_),
    .Q(net354),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43813_ (.D(_03657_),
    .Q(net355),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_4 _43814_ (.D(_03658_),
    .Q(net356),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_4 _43815_ (.D(_03659_),
    .Q(net357),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_4 _43816_ (.D(_03660_),
    .Q(net358),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_4 _43817_ (.D(_03661_),
    .Q(net359),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_4 _43818_ (.D(_03662_),
    .Q(net361),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_4 _43819_ (.D(_03663_),
    .Q(net362),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 _43820_ (.D(_03664_),
    .Q(\cpuregs[9][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43821_ (.D(_03665_),
    .Q(\cpuregs[9][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43822_ (.D(_03666_),
    .Q(\cpuregs[9][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43823_ (.D(_03667_),
    .Q(\cpuregs[9][3] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43824_ (.D(_03668_),
    .Q(\cpuregs[9][4] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43825_ (.D(_03669_),
    .Q(\cpuregs[9][5] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43826_ (.D(_03670_),
    .Q(\cpuregs[9][6] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43827_ (.D(_03671_),
    .Q(\cpuregs[9][7] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43828_ (.D(_03672_),
    .Q(\cpuregs[9][8] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43829_ (.D(_03673_),
    .Q(\cpuregs[9][9] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43830_ (.D(_03674_),
    .Q(\cpuregs[9][10] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43831_ (.D(_03675_),
    .Q(\cpuregs[9][11] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43832_ (.D(_03676_),
    .Q(\cpuregs[9][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43833_ (.D(_03677_),
    .Q(\cpuregs[9][13] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _43834_ (.D(_03678_),
    .Q(\cpuregs[9][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43835_ (.D(_03679_),
    .Q(\cpuregs[9][15] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43836_ (.D(_03680_),
    .Q(\cpuregs[9][16] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _43837_ (.D(_03681_),
    .Q(\cpuregs[9][17] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_1 _43838_ (.D(_03682_),
    .Q(\cpuregs[9][18] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__dfxtp_1 _43839_ (.D(_03683_),
    .Q(\cpuregs[9][19] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__dfxtp_1 _43840_ (.D(_03684_),
    .Q(\cpuregs[9][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43841_ (.D(_03685_),
    .Q(\cpuregs[9][21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43842_ (.D(_03686_),
    .Q(\cpuregs[9][22] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _43843_ (.D(_03687_),
    .Q(\cpuregs[9][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43844_ (.D(_03688_),
    .Q(\cpuregs[9][24] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 _43845_ (.D(_03689_),
    .Q(\cpuregs[9][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43846_ (.D(_03690_),
    .Q(\cpuregs[9][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43847_ (.D(_03691_),
    .Q(\cpuregs[9][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43848_ (.D(_03692_),
    .Q(\cpuregs[9][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43849_ (.D(_03693_),
    .Q(\cpuregs[9][29] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43850_ (.D(_03694_),
    .Q(\cpuregs[9][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43851_ (.D(_03695_),
    .Q(\cpuregs[9][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43852_ (.D(_03696_),
    .Q(\cpuregs[6][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43853_ (.D(_03697_),
    .Q(\cpuregs[6][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _43854_ (.D(_03698_),
    .Q(\cpuregs[6][2] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43855_ (.D(_03699_),
    .Q(\cpuregs[6][3] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43856_ (.D(_03700_),
    .Q(\cpuregs[6][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43857_ (.D(_03701_),
    .Q(\cpuregs[6][5] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43858_ (.D(_03702_),
    .Q(\cpuregs[6][6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43859_ (.D(_03703_),
    .Q(\cpuregs[6][7] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43860_ (.D(_03704_),
    .Q(\cpuregs[6][8] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43861_ (.D(_03705_),
    .Q(\cpuregs[6][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43862_ (.D(_03706_),
    .Q(\cpuregs[6][10] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43863_ (.D(_03707_),
    .Q(\cpuregs[6][11] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43864_ (.D(_03708_),
    .Q(\cpuregs[6][12] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43865_ (.D(_03709_),
    .Q(\cpuregs[6][13] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43866_ (.D(_03710_),
    .Q(\cpuregs[6][14] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43867_ (.D(_03711_),
    .Q(\cpuregs[6][15] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43868_ (.D(_03712_),
    .Q(\cpuregs[6][16] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_1 _43869_ (.D(_03713_),
    .Q(\cpuregs[6][17] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43870_ (.D(_03714_),
    .Q(\cpuregs[6][18] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43871_ (.D(_03715_),
    .Q(\cpuregs[6][19] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__dfxtp_1 _43872_ (.D(_03716_),
    .Q(\cpuregs[6][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43873_ (.D(_03717_),
    .Q(\cpuregs[6][21] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43874_ (.D(_03718_),
    .Q(\cpuregs[6][22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _43875_ (.D(_03719_),
    .Q(\cpuregs[6][23] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43876_ (.D(_03720_),
    .Q(\cpuregs[6][24] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _43877_ (.D(_03721_),
    .Q(\cpuregs[6][25] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _43878_ (.D(_03722_),
    .Q(\cpuregs[6][26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43879_ (.D(_03723_),
    .Q(\cpuregs[6][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43880_ (.D(_03724_),
    .Q(\cpuregs[6][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43881_ (.D(_03725_),
    .Q(\cpuregs[6][29] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43882_ (.D(_03726_),
    .Q(\cpuregs[6][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43883_ (.D(_03727_),
    .Q(\cpuregs[6][31] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43884_ (.D(_03728_),
    .Q(\pcpi_mul.active[0] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_2 _43885_ (.D(_03729_),
    .Q(\pcpi_mul.active[1] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_4 _43886_ (.D(_03730_),
    .Q(net408),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_2 _43887_ (.D(_03731_),
    .Q(\count_cycle[0] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43888_ (.D(_03732_),
    .Q(\count_cycle[1] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43889_ (.D(_03733_),
    .Q(\count_cycle[2] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43890_ (.D(_03734_),
    .Q(\count_cycle[3] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43891_ (.D(_03735_),
    .Q(\count_cycle[4] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43892_ (.D(_03736_),
    .Q(\count_cycle[5] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43893_ (.D(_03737_),
    .Q(\count_cycle[6] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43894_ (.D(_03738_),
    .Q(\count_cycle[7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43895_ (.D(_03739_),
    .Q(\count_cycle[8] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43896_ (.D(_03740_),
    .Q(\count_cycle[9] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43897_ (.D(_03741_),
    .Q(\count_cycle[10] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43898_ (.D(_03742_),
    .Q(\count_cycle[11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43899_ (.D(_03743_),
    .Q(\count_cycle[12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43900_ (.D(_03744_),
    .Q(\count_cycle[13] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43901_ (.D(_03745_),
    .Q(\count_cycle[14] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43902_ (.D(_03746_),
    .Q(\count_cycle[15] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43903_ (.D(_03747_),
    .Q(\count_cycle[16] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43904_ (.D(_03748_),
    .Q(\count_cycle[17] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43905_ (.D(_03749_),
    .Q(\count_cycle[18] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43906_ (.D(_03750_),
    .Q(\count_cycle[19] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43907_ (.D(_03751_),
    .Q(\count_cycle[20] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43908_ (.D(_03752_),
    .Q(\count_cycle[21] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43909_ (.D(_03753_),
    .Q(\count_cycle[22] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _43910_ (.D(_03754_),
    .Q(\count_cycle[23] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _43911_ (.D(_03755_),
    .Q(\count_cycle[24] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43912_ (.D(_03756_),
    .Q(\count_cycle[25] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43913_ (.D(_03757_),
    .Q(\count_cycle[26] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43914_ (.D(_03758_),
    .Q(\count_cycle[27] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43915_ (.D(_03759_),
    .Q(\count_cycle[28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43916_ (.D(_03760_),
    .Q(\count_cycle[29] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43917_ (.D(_03761_),
    .Q(\count_cycle[30] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43918_ (.D(_03762_),
    .Q(\count_cycle[31] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43919_ (.D(_03763_),
    .Q(\count_cycle[32] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43920_ (.D(_03764_),
    .Q(\count_cycle[33] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43921_ (.D(_03765_),
    .Q(\count_cycle[34] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43922_ (.D(_03766_),
    .Q(\count_cycle[35] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43923_ (.D(_03767_),
    .Q(\count_cycle[36] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43924_ (.D(_03768_),
    .Q(\count_cycle[37] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43925_ (.D(_03769_),
    .Q(\count_cycle[38] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43926_ (.D(_03770_),
    .Q(\count_cycle[39] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43927_ (.D(_03771_),
    .Q(\count_cycle[40] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43928_ (.D(_03772_),
    .Q(\count_cycle[41] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43929_ (.D(_03773_),
    .Q(\count_cycle[42] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43930_ (.D(_03774_),
    .Q(\count_cycle[43] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43931_ (.D(_03775_),
    .Q(\count_cycle[44] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43932_ (.D(_03776_),
    .Q(\count_cycle[45] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _43933_ (.D(_03777_),
    .Q(\count_cycle[46] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _43934_ (.D(_03778_),
    .Q(\count_cycle[47] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _43935_ (.D(_03779_),
    .Q(\count_cycle[48] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _43936_ (.D(_03780_),
    .Q(\count_cycle[49] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _43937_ (.D(_03781_),
    .Q(\count_cycle[50] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _43938_ (.D(_03782_),
    .Q(\count_cycle[51] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _43939_ (.D(_03783_),
    .Q(\count_cycle[52] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _43940_ (.D(_03784_),
    .Q(\count_cycle[53] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _43941_ (.D(_03785_),
    .Q(\count_cycle[54] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _43942_ (.D(_03786_),
    .Q(\count_cycle[55] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _43943_ (.D(_03787_),
    .Q(\count_cycle[56] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 _43944_ (.D(_03788_),
    .Q(\count_cycle[57] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _43945_ (.D(_03789_),
    .Q(\count_cycle[58] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _43946_ (.D(_03790_),
    .Q(\count_cycle[59] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43947_ (.D(_03791_),
    .Q(\count_cycle[60] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _43948_ (.D(_03792_),
    .Q(\count_cycle[61] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _43949_ (.D(_03793_),
    .Q(\count_cycle[62] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 _43950_ (.D(_03794_),
    .Q(\count_cycle[63] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _43951_ (.D(_03795_),
    .Q(\timer[0] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43952_ (.D(_03796_),
    .Q(\timer[1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43953_ (.D(_03797_),
    .Q(\timer[2] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _43954_ (.D(_03798_),
    .Q(\timer[3] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43955_ (.D(_03799_),
    .Q(\timer[4] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43956_ (.D(_03800_),
    .Q(\timer[5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43957_ (.D(_03801_),
    .Q(\timer[6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43958_ (.D(_03802_),
    .Q(\timer[7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43959_ (.D(_03803_),
    .Q(\timer[8] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43960_ (.D(_03804_),
    .Q(\timer[9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43961_ (.D(_03805_),
    .Q(\timer[10] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43962_ (.D(_03806_),
    .Q(\timer[11] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43963_ (.D(_03807_),
    .Q(\timer[12] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43964_ (.D(_03808_),
    .Q(\timer[13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43965_ (.D(_03809_),
    .Q(\timer[14] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43966_ (.D(_03810_),
    .Q(\timer[15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43967_ (.D(_03811_),
    .Q(\timer[16] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43968_ (.D(_03812_),
    .Q(\timer[17] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43969_ (.D(_03813_),
    .Q(\timer[18] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43970_ (.D(_03814_),
    .Q(\timer[19] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43971_ (.D(_03815_),
    .Q(\timer[20] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43972_ (.D(_03816_),
    .Q(\timer[21] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43973_ (.D(_03817_),
    .Q(\timer[22] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43974_ (.D(_03818_),
    .Q(\timer[23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43975_ (.D(_03819_),
    .Q(\timer[24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43976_ (.D(_03820_),
    .Q(\timer[25] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43977_ (.D(_03821_),
    .Q(\timer[26] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _43978_ (.D(_03822_),
    .Q(\timer[27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43979_ (.D(_03823_),
    .Q(\timer[28] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43980_ (.D(_03824_),
    .Q(\timer[29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43981_ (.D(_03825_),
    .Q(\timer[30] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43982_ (.D(_03826_),
    .Q(\timer[31] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43983_ (.D(_03827_),
    .Q(pcpi_timeout),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _43984_ (.D(_03828_),
    .Q(decoder_pseudo_trigger),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_2 _43985_ (.D(_03829_),
    .Q(is_compare),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 _43986_ (.D(_03830_),
    .Q(do_waitirq),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_4 _43987_ (.D(_03831_),
    .Q(net237),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_4 _43988_ (.D(_03832_),
    .Q(net370),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_4 _43989_ (.D(_03833_),
    .Q(net102),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_4 _43990_ (.D(_03834_),
    .Q(net113),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 _43991_ (.D(_03835_),
    .Q(net124),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _43992_ (.D(_03836_),
    .Q(net127),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _43993_ (.D(_03837_),
    .Q(net128),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _43994_ (.D(_03838_),
    .Q(net129),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_4 _43995_ (.D(_03839_),
    .Q(net130),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _43996_ (.D(_03840_),
    .Q(net131),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _43997_ (.D(_03841_),
    .Q(net132),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 _43998_ (.D(_03842_),
    .Q(net133),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _43999_ (.D(_03843_),
    .Q(net103),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _44000_ (.D(_03844_),
    .Q(net104),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 _44001_ (.D(_03845_),
    .Q(net105),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _44002_ (.D(_03846_),
    .Q(net106),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _44003_ (.D(_03847_),
    .Q(net107),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 _44004_ (.D(_03848_),
    .Q(net108),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _44005_ (.D(_03849_),
    .Q(net109),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_4 _44006_ (.D(_03850_),
    .Q(net110),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _44007_ (.D(_03851_),
    .Q(net111),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _44008_ (.D(_03852_),
    .Q(net112),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_4 _44009_ (.D(_03853_),
    .Q(net114),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_4 _44010_ (.D(_03854_),
    .Q(net115),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _44011_ (.D(_03855_),
    .Q(net116),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_4 _44012_ (.D(_03856_),
    .Q(net117),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_2 _44013_ (.D(_03857_),
    .Q(net118),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _44014_ (.D(_03858_),
    .Q(net119),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_4 _44015_ (.D(_03859_),
    .Q(net120),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_4 _44016_ (.D(_03860_),
    .Q(net121),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_4 _44017_ (.D(_03861_),
    .Q(net122),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_4 _44018_ (.D(_03862_),
    .Q(net123),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _44019_ (.D(_03863_),
    .Q(net125),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_4 _44020_ (.D(_03864_),
    .Q(net126),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _44021_ (.D(_03865_),
    .Q(\count_instr[0] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _44022_ (.D(_03866_),
    .Q(\count_instr[1] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _44023_ (.D(_03867_),
    .Q(\count_instr[2] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _44024_ (.D(_03868_),
    .Q(\count_instr[3] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _44025_ (.D(_03869_),
    .Q(\count_instr[4] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _44026_ (.D(_03870_),
    .Q(\count_instr[5] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _44027_ (.D(_03871_),
    .Q(\count_instr[6] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _44028_ (.D(_03872_),
    .Q(\count_instr[7] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _44029_ (.D(_03873_),
    .Q(\count_instr[8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _44030_ (.D(_03874_),
    .Q(\count_instr[9] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _44031_ (.D(_03875_),
    .Q(\count_instr[10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _44032_ (.D(_03876_),
    .Q(\count_instr[11] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _44033_ (.D(_03877_),
    .Q(\count_instr[12] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44034_ (.D(_03878_),
    .Q(\count_instr[13] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44035_ (.D(_03879_),
    .Q(\count_instr[14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _44036_ (.D(_03880_),
    .Q(\count_instr[15] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _44037_ (.D(_03881_),
    .Q(\count_instr[16] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _44038_ (.D(_03882_),
    .Q(\count_instr[17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _44039_ (.D(_03883_),
    .Q(\count_instr[18] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44040_ (.D(_03884_),
    .Q(\count_instr[19] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44041_ (.D(_03885_),
    .Q(\count_instr[20] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44042_ (.D(_03886_),
    .Q(\count_instr[21] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44043_ (.D(_03887_),
    .Q(\count_instr[22] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44044_ (.D(_03888_),
    .Q(\count_instr[23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44045_ (.D(_03889_),
    .Q(\count_instr[24] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44046_ (.D(_03890_),
    .Q(\count_instr[25] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44047_ (.D(_03891_),
    .Q(\count_instr[26] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44048_ (.D(_03892_),
    .Q(\count_instr[27] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44049_ (.D(_03893_),
    .Q(\count_instr[28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44050_ (.D(_03894_),
    .Q(\count_instr[29] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44051_ (.D(_03895_),
    .Q(\count_instr[30] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _44052_ (.D(_03896_),
    .Q(\count_instr[31] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _44053_ (.D(_03897_),
    .Q(\count_instr[32] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44054_ (.D(_03898_),
    .Q(\count_instr[33] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44055_ (.D(_03899_),
    .Q(\count_instr[34] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44056_ (.D(_03900_),
    .Q(\count_instr[35] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _44057_ (.D(_03901_),
    .Q(\count_instr[36] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44058_ (.D(_03902_),
    .Q(\count_instr[37] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _44059_ (.D(_03903_),
    .Q(\count_instr[38] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _44060_ (.D(_03904_),
    .Q(\count_instr[39] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _44061_ (.D(_03905_),
    .Q(\count_instr[40] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44062_ (.D(_03906_),
    .Q(\count_instr[41] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44063_ (.D(_03907_),
    .Q(\count_instr[42] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44064_ (.D(_03908_),
    .Q(\count_instr[43] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _44065_ (.D(_03909_),
    .Q(\count_instr[44] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _44066_ (.D(_03910_),
    .Q(\count_instr[45] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 _44067_ (.D(_03911_),
    .Q(\count_instr[46] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _44068_ (.D(_03912_),
    .Q(\count_instr[47] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 _44069_ (.D(_03913_),
    .Q(\count_instr[48] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _44070_ (.D(_03914_),
    .Q(\count_instr[49] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_2 _44071_ (.D(_03915_),
    .Q(\count_instr[50] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _44072_ (.D(_03916_),
    .Q(\count_instr[51] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _44073_ (.D(_03917_),
    .Q(\count_instr[52] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44074_ (.D(_03918_),
    .Q(\count_instr[53] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _44075_ (.D(_03919_),
    .Q(\count_instr[54] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 _44076_ (.D(_03920_),
    .Q(\count_instr[55] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44077_ (.D(_03921_),
    .Q(\count_instr[56] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 _44078_ (.D(_03922_),
    .Q(\count_instr[57] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 _44079_ (.D(_03923_),
    .Q(\count_instr[58] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44080_ (.D(_03924_),
    .Q(\count_instr[59] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44081_ (.D(_03925_),
    .Q(\count_instr[60] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44082_ (.D(_03926_),
    .Q(\count_instr[61] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 _44083_ (.D(_03927_),
    .Q(\count_instr[62] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 _44084_ (.D(_03928_),
    .Q(\count_instr[63] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _44085_ (.D(_03929_),
    .Q(\reg_pc[1] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 _44086_ (.D(_03930_),
    .Q(\reg_pc[2] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 _44087_ (.D(_03931_),
    .Q(\reg_pc[3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _44088_ (.D(_03932_),
    .Q(\reg_pc[4] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _44089_ (.D(_03933_),
    .Q(\reg_pc[5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _44090_ (.D(_03934_),
    .Q(\reg_pc[6] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _44091_ (.D(_03935_),
    .Q(\reg_pc[7] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _44092_ (.D(_03936_),
    .Q(\reg_pc[8] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _44093_ (.D(_03937_),
    .Q(\reg_pc[9] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _44094_ (.D(_03938_),
    .Q(\reg_pc[10] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _44095_ (.D(_03939_),
    .Q(\reg_pc[11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _44096_ (.D(_03940_),
    .Q(\reg_pc[12] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _44097_ (.D(_03941_),
    .Q(\reg_pc[13] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _44098_ (.D(_03942_),
    .Q(\reg_pc[14] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _44099_ (.D(_03943_),
    .Q(\reg_pc[15] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 _44100_ (.D(_03944_),
    .Q(\reg_pc[16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_2 _44101_ (.D(_03945_),
    .Q(\reg_pc[17] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _44102_ (.D(_03946_),
    .Q(\reg_pc[18] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _44103_ (.D(_03947_),
    .Q(\reg_pc[19] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _44104_ (.D(_03948_),
    .Q(\reg_pc[20] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _44105_ (.D(_03949_),
    .Q(\reg_pc[21] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _44106_ (.D(_03950_),
    .Q(\reg_pc[22] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _44107_ (.D(_03951_),
    .Q(\reg_pc[23] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _44108_ (.D(_03952_),
    .Q(\reg_pc[24] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _44109_ (.D(_03953_),
    .Q(\reg_pc[25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _44110_ (.D(_03954_),
    .Q(\reg_pc[26] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _44111_ (.D(_03955_),
    .Q(\reg_pc[27] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _44112_ (.D(_03956_),
    .Q(\reg_pc[28] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _44113_ (.D(_03957_),
    .Q(\reg_pc[29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _44114_ (.D(_03958_),
    .Q(\reg_pc[30] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _44115_ (.D(_03959_),
    .Q(\reg_pc[31] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _44116_ (.D(_03960_),
    .Q(\reg_next_pc[1] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 _44117_ (.D(_03961_),
    .Q(\reg_next_pc[2] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 _44118_ (.D(_03962_),
    .Q(\reg_next_pc[3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _44119_ (.D(_03963_),
    .Q(\reg_next_pc[4] ),
    .CLK(clknet_5_18_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _44120_ (.D(_03964_),
    .Q(\reg_next_pc[5] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _44121_ (.D(_03965_),
    .Q(\reg_next_pc[6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 _44122_ (.D(_03966_),
    .Q(\reg_next_pc[7] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _44123_ (.D(_03967_),
    .Q(\reg_next_pc[8] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _44124_ (.D(_03968_),
    .Q(\reg_next_pc[9] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _44125_ (.D(_03969_),
    .Q(\reg_next_pc[10] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _44126_ (.D(_03970_),
    .Q(\reg_next_pc[11] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _44127_ (.D(_03971_),
    .Q(\reg_next_pc[12] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _44128_ (.D(_03972_),
    .Q(\reg_next_pc[13] ),
    .CLK(clknet_5_18_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _44129_ (.D(_03973_),
    .Q(\reg_next_pc[14] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_1 _44130_ (.D(_03974_),
    .Q(\reg_next_pc[15] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _44131_ (.D(_03975_),
    .Q(\reg_next_pc[16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _44132_ (.D(_03976_),
    .Q(\reg_next_pc[17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _44133_ (.D(_03977_),
    .Q(\reg_next_pc[18] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _44134_ (.D(_03978_),
    .Q(\reg_next_pc[19] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_1 _44135_ (.D(_03979_),
    .Q(\reg_next_pc[20] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_1 _44136_ (.D(_03980_),
    .Q(\reg_next_pc[21] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_1 _44137_ (.D(_03981_),
    .Q(\reg_next_pc[22] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _44138_ (.D(_03982_),
    .Q(\reg_next_pc[23] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _44139_ (.D(_03983_),
    .Q(\reg_next_pc[24] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _44140_ (.D(_03984_),
    .Q(\reg_next_pc[25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _44141_ (.D(_03985_),
    .Q(\reg_next_pc[26] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _44142_ (.D(_03986_),
    .Q(\reg_next_pc[27] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _44143_ (.D(_03987_),
    .Q(\reg_next_pc[28] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _44144_ (.D(_03988_),
    .Q(\reg_next_pc[29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _44145_ (.D(_03989_),
    .Q(\reg_next_pc[30] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _44146_ (.D(_03990_),
    .Q(\reg_next_pc[31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _44147_ (.D(_03991_),
    .Q(mem_do_rdata),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _44148_ (.D(_03992_),
    .Q(mem_do_wdata),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _44149_ (.D(_03993_),
    .Q(\pcpi_timeout_counter[0] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _44150_ (.D(_03994_),
    .Q(\pcpi_timeout_counter[1] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _44151_ (.D(_03995_),
    .Q(\pcpi_timeout_counter[2] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 _44152_ (.D(_03996_),
    .Q(\pcpi_timeout_counter[3] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 _44153_ (.D(_03997_),
    .Q(instr_beq),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _44154_ (.D(_03998_),
    .Q(instr_bne),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _44155_ (.D(_03999_),
    .Q(instr_blt),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _44156_ (.D(_04000_),
    .Q(instr_bge),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _44157_ (.D(_04001_),
    .Q(instr_bltu),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _44158_ (.D(_04002_),
    .Q(instr_bgeu),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _44159_ (.D(_04003_),
    .Q(instr_addi),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _44160_ (.D(_04004_),
    .Q(instr_slti),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _44161_ (.D(_04005_),
    .Q(instr_sltiu),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _44162_ (.D(_04006_),
    .Q(instr_xori),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_2 _44163_ (.D(_04007_),
    .Q(instr_ori),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _44164_ (.D(_04008_),
    .Q(instr_andi),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _44165_ (.D(_04009_),
    .Q(instr_add),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_4 _44166_ (.D(_04010_),
    .Q(instr_sub),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _44167_ (.D(_04011_),
    .Q(instr_sll),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _44168_ (.D(_04012_),
    .Q(instr_slt),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_1 _44169_ (.D(_04013_),
    .Q(instr_sltu),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _44170_ (.D(_04014_),
    .Q(instr_xor),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _44171_ (.D(_04015_),
    .Q(instr_srl),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _44172_ (.D(_04016_),
    .Q(instr_sra),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _44173_ (.D(_04017_),
    .Q(instr_or),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _44174_ (.D(_04018_),
    .Q(instr_and),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _44175_ (.D(_04019_),
    .Q(\decoded_rs1[0] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 _44176_ (.D(_04020_),
    .Q(\decoded_rs1[1] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 _44177_ (.D(_04021_),
    .Q(\decoded_rs1[2] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 _44178_ (.D(_04022_),
    .Q(\decoded_rs1[3] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 _44179_ (.D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 _44180_ (.D(_04024_),
    .Q(net166),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _44181_ (.D(_04025_),
    .Q(\irq_mask[0] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _44182_ (.D(_04026_),
    .Q(\irq_mask[1] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _44183_ (.D(_04027_),
    .Q(\irq_mask[2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _44184_ (.D(_04028_),
    .Q(\irq_mask[3] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _44185_ (.D(_04029_),
    .Q(\irq_mask[4] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _44186_ (.D(_04030_),
    .Q(\irq_mask[5] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _44187_ (.D(_04031_),
    .Q(\irq_mask[6] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _44188_ (.D(_04032_),
    .Q(\irq_mask[7] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _44189_ (.D(_04033_),
    .Q(\irq_mask[8] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _44190_ (.D(_04034_),
    .Q(\irq_mask[9] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _44191_ (.D(_04035_),
    .Q(\irq_mask[10] ),
    .CLK(clknet_5_16_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _44192_ (.D(_04036_),
    .Q(\irq_mask[11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _44193_ (.D(_04037_),
    .Q(\irq_mask[12] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _44194_ (.D(_04038_),
    .Q(\irq_mask[13] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _44195_ (.D(_04039_),
    .Q(\irq_mask[14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _44196_ (.D(_04040_),
    .Q(\irq_mask[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _44197_ (.D(_04041_),
    .Q(\irq_mask[16] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _44198_ (.D(_04042_),
    .Q(\irq_mask[17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _44199_ (.D(_04043_),
    .Q(\irq_mask[18] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _44200_ (.D(_04044_),
    .Q(\irq_mask[19] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _44201_ (.D(_04045_),
    .Q(\irq_mask[20] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _44202_ (.D(_04046_),
    .Q(\irq_mask[21] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _44203_ (.D(_04047_),
    .Q(\irq_mask[22] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _44204_ (.D(_04048_),
    .Q(\irq_mask[23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _44205_ (.D(_04049_),
    .Q(\irq_mask[24] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _44206_ (.D(_04050_),
    .Q(\irq_mask[25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _44207_ (.D(_04051_),
    .Q(\irq_mask[26] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _44208_ (.D(_04052_),
    .Q(\irq_mask[27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _44209_ (.D(_04053_),
    .Q(\irq_mask[28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _44210_ (.D(_04054_),
    .Q(\irq_mask[29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _44211_ (.D(_04055_),
    .Q(\irq_mask[30] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _44212_ (.D(_04056_),
    .Q(\irq_mask[31] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _44213_ (.D(_04057_),
    .Q(mem_do_prefetch),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _44214_ (.D(_04058_),
    .Q(mem_do_rinst),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _44215_ (.D(_04059_),
    .Q(\irq_state[0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _44216_ (.D(_04060_),
    .Q(\irq_state[1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _44217_ (.D(_04061_),
    .Q(latched_store),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_4 _44218_ (.D(_04062_),
    .Q(latched_stalu),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_4 _44219_ (.D(_04063_),
    .Q(\pcpi_mul.rs2[32] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _44220_ (.D(_04064_),
    .Q(\pcpi_mul.rs1[32] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 _44221_ (.D(_04065_),
    .Q(irq_delay),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _44222_ (.D(_04066_),
    .Q(\decoded_rs1[4] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_2 _44223_ (.D(_04067_),
    .Q(\mem_state[0] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_2 _44224_ (.D(_04068_),
    .Q(\mem_state[1] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_4 _44225_ (.D(_04069_),
    .Q(latched_branch),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _44226_ (.D(_04070_),
    .Q(latched_is_lh),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _44227_ (.D(_04071_),
    .Q(latched_is_lb),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _44228_ (.D(_04072_),
    .Q(irq_active),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8859 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(irq[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(irq[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(irq[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(irq[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(irq[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(irq[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(irq[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(irq[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(irq[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(irq[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(irq[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(irq[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(irq[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_8 input14 (.A(irq[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(irq[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(irq[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(irq[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(irq[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(irq[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(irq[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(irq[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input22 (.A(irq[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(irq[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_6 input24 (.A(irq[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_8 input25 (.A(irq[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(irq[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_8 input27 (.A(irq[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(irq[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_8 input29 (.A(irq[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(irq[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(irq[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_6 input32 (.A(irq[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(mem_rdata[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(mem_rdata[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(mem_rdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(mem_rdata[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(mem_rdata[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(mem_rdata[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(mem_rdata[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input40 (.A(mem_rdata[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_6 input41 (.A(mem_rdata[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(mem_rdata[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(mem_rdata[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(mem_rdata[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(mem_rdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(mem_rdata[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_8 input47 (.A(mem_rdata[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(mem_rdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(mem_rdata[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_8 input50 (.A(mem_rdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(mem_rdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(mem_rdata[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_6 input53 (.A(mem_rdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_8 input54 (.A(mem_rdata[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 input55 (.A(mem_rdata[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(mem_rdata[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_8 input57 (.A(mem_rdata[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input58 (.A(mem_rdata[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(mem_rdata[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(mem_rdata[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(mem_rdata[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(mem_rdata[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(mem_rdata[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(mem_rdata[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(mem_ready),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(pcpi_rd[0]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(pcpi_rd[10]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(pcpi_rd[11]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(pcpi_rd[12]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(pcpi_rd[13]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(pcpi_rd[14]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(pcpi_rd[15]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(pcpi_rd[16]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(pcpi_rd[17]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(pcpi_rd[18]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(pcpi_rd[19]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(pcpi_rd[1]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(pcpi_rd[20]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(pcpi_rd[21]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(pcpi_rd[22]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(pcpi_rd[23]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(pcpi_rd[24]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(pcpi_rd[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(pcpi_rd[26]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(pcpi_rd[27]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(pcpi_rd[28]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(pcpi_rd[29]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(pcpi_rd[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(pcpi_rd[30]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(pcpi_rd[31]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(pcpi_rd[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(pcpi_rd[4]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(pcpi_rd[5]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(pcpi_rd[6]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(pcpi_rd[7]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(pcpi_rd[8]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(pcpi_rd[9]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(pcpi_ready),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(pcpi_wait),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(pcpi_wr),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 input101 (.A(resetn),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(eoi[0]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(eoi[10]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(eoi[11]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(eoi[12]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(eoi[13]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(eoi[14]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(eoi[15]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(eoi[16]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(eoi[17]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(eoi[18]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(eoi[19]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(eoi[1]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(eoi[20]));
 sky130_fd_sc_hd__clkbuf_2 output115 (.A(net115),
    .X(eoi[21]));
 sky130_fd_sc_hd__clkbuf_2 output116 (.A(net116),
    .X(eoi[22]));
 sky130_fd_sc_hd__clkbuf_2 output117 (.A(net117),
    .X(eoi[23]));
 sky130_fd_sc_hd__clkbuf_2 output118 (.A(net118),
    .X(eoi[24]));
 sky130_fd_sc_hd__clkbuf_2 output119 (.A(net119),
    .X(eoi[25]));
 sky130_fd_sc_hd__clkbuf_2 output120 (.A(net120),
    .X(eoi[26]));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(eoi[27]));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(eoi[28]));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(eoi[29]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(eoi[2]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(eoi[30]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(eoi[31]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(eoi[3]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(eoi[4]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(eoi[5]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(eoi[6]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(eoi[7]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(eoi[8]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(eoi[9]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output161 (.A(net161),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output162 (.A(net162),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output163 (.A(net163),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output164 (.A(net164),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output165 (.A(net165),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output166 (.A(net166),
    .X(mem_instr));
 sky130_fd_sc_hd__clkbuf_2 output167 (.A(net167),
    .X(mem_la_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output168 (.A(net168),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output169 (.A(net169),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output170 (.A(net170),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output171 (.A(net171),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output172 (.A(net172),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output173 (.A(net173),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output174 (.A(net174),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output175 (.A(net175),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output176 (.A(net176),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output177 (.A(net177),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output178 (.A(net178),
    .X(mem_la_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output179 (.A(net179),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output180 (.A(net180),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output181 (.A(net181),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output182 (.A(net182),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output183 (.A(net183),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output184 (.A(net184),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output185 (.A(net185),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output186 (.A(net186),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output187 (.A(net187),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output188 (.A(net188),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output189 (.A(net189),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output190 (.A(net190),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output191 (.A(net191),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output192 (.A(net192),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output193 (.A(net193),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output194 (.A(net194),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output195 (.A(net195),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output196 (.A(net196),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output197 (.A(net197),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output198 (.A(net198),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output199 (.A(net199),
    .X(mem_la_read));
 sky130_fd_sc_hd__clkbuf_2 output200 (.A(net516),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output201 (.A(net201),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output202 (.A(net202),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output203 (.A(net203),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output204 (.A(net204),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output205 (.A(net205),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output215 (.A(net215),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output216 (.A(net216),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output217 (.A(net217),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output218 (.A(net435),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net514),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output223 (.A(net223),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output224 (.A(net224),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output225 (.A(net225),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output226 (.A(net226),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output227 (.A(net227),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output228 (.A(net228),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output229 (.A(net229),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output232 (.A(net232),
    .X(mem_la_write));
 sky130_fd_sc_hd__clkbuf_2 output233 (.A(net233),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output234 (.A(net234),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net235),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output236 (.A(net236),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output237 (.A(net237),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_2 output238 (.A(net238),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output239 (.A(net239),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output240 (.A(net240),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output241 (.A(net241),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output242 (.A(net242),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output243 (.A(net243),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output244 (.A(net244),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output245 (.A(net245),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output246 (.A(net246),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output247 (.A(net247),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output248 (.A(net248),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output249 (.A(net249),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output250 (.A(net250),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output251 (.A(net251),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output252 (.A(net252),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output253 (.A(net253),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output254 (.A(net254),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output255 (.A(net255),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output256 (.A(net256),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output257 (.A(net257),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output258 (.A(net258),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output259 (.A(net259),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output260 (.A(net260),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output261 (.A(net261),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output262 (.A(net262),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output263 (.A(net263),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output265 (.A(net265),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output266 (.A(net266),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output267 (.A(net267),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output268 (.A(net268),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output269 (.A(net269),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output271 (.A(net271),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output272 (.A(net272),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output273 (.A(net273),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output274 (.A(net274),
    .X(pcpi_insn[0]));
 sky130_fd_sc_hd__clkbuf_2 output275 (.A(net275),
    .X(pcpi_insn[10]));
 sky130_fd_sc_hd__clkbuf_2 output276 (.A(net276),
    .X(pcpi_insn[11]));
 sky130_fd_sc_hd__clkbuf_2 output277 (.A(net277),
    .X(pcpi_insn[12]));
 sky130_fd_sc_hd__clkbuf_2 output278 (.A(net278),
    .X(pcpi_insn[13]));
 sky130_fd_sc_hd__clkbuf_2 output279 (.A(net279),
    .X(pcpi_insn[14]));
 sky130_fd_sc_hd__clkbuf_2 output280 (.A(net280),
    .X(pcpi_insn[15]));
 sky130_fd_sc_hd__clkbuf_2 output281 (.A(net281),
    .X(pcpi_insn[16]));
 sky130_fd_sc_hd__clkbuf_2 output282 (.A(net282),
    .X(pcpi_insn[17]));
 sky130_fd_sc_hd__clkbuf_2 output283 (.A(net283),
    .X(pcpi_insn[18]));
 sky130_fd_sc_hd__clkbuf_2 output284 (.A(net284),
    .X(pcpi_insn[19]));
 sky130_fd_sc_hd__clkbuf_2 output285 (.A(net285),
    .X(pcpi_insn[1]));
 sky130_fd_sc_hd__clkbuf_2 output286 (.A(net286),
    .X(pcpi_insn[20]));
 sky130_fd_sc_hd__clkbuf_2 output287 (.A(net287),
    .X(pcpi_insn[21]));
 sky130_fd_sc_hd__clkbuf_2 output288 (.A(net288),
    .X(pcpi_insn[22]));
 sky130_fd_sc_hd__clkbuf_2 output289 (.A(net289),
    .X(pcpi_insn[23]));
 sky130_fd_sc_hd__clkbuf_2 output290 (.A(net290),
    .X(pcpi_insn[24]));
 sky130_fd_sc_hd__clkbuf_2 output291 (.A(net291),
    .X(pcpi_insn[25]));
 sky130_fd_sc_hd__clkbuf_2 output292 (.A(net292),
    .X(pcpi_insn[26]));
 sky130_fd_sc_hd__clkbuf_2 output293 (.A(net293),
    .X(pcpi_insn[27]));
 sky130_fd_sc_hd__clkbuf_2 output294 (.A(net294),
    .X(pcpi_insn[28]));
 sky130_fd_sc_hd__clkbuf_2 output295 (.A(net295),
    .X(pcpi_insn[29]));
 sky130_fd_sc_hd__clkbuf_2 output296 (.A(net296),
    .X(pcpi_insn[2]));
 sky130_fd_sc_hd__clkbuf_2 output297 (.A(net297),
    .X(pcpi_insn[30]));
 sky130_fd_sc_hd__clkbuf_2 output298 (.A(net298),
    .X(pcpi_insn[31]));
 sky130_fd_sc_hd__clkbuf_2 output299 (.A(net299),
    .X(pcpi_insn[3]));
 sky130_fd_sc_hd__clkbuf_2 output300 (.A(net300),
    .X(pcpi_insn[4]));
 sky130_fd_sc_hd__clkbuf_2 output301 (.A(net301),
    .X(pcpi_insn[5]));
 sky130_fd_sc_hd__clkbuf_2 output302 (.A(net302),
    .X(pcpi_insn[6]));
 sky130_fd_sc_hd__clkbuf_2 output303 (.A(net303),
    .X(pcpi_insn[7]));
 sky130_fd_sc_hd__clkbuf_2 output304 (.A(net304),
    .X(pcpi_insn[8]));
 sky130_fd_sc_hd__clkbuf_2 output305 (.A(net305),
    .X(pcpi_insn[9]));
 sky130_fd_sc_hd__clkbuf_2 output306 (.A(net306),
    .X(pcpi_rs1[0]));
 sky130_fd_sc_hd__clkbuf_2 output307 (.A(net307),
    .X(pcpi_rs1[10]));
 sky130_fd_sc_hd__clkbuf_2 output308 (.A(net308),
    .X(pcpi_rs1[11]));
 sky130_fd_sc_hd__clkbuf_2 output309 (.A(net309),
    .X(pcpi_rs1[12]));
 sky130_fd_sc_hd__clkbuf_2 output310 (.A(net310),
    .X(pcpi_rs1[13]));
 sky130_fd_sc_hd__clkbuf_2 output311 (.A(net311),
    .X(pcpi_rs1[14]));
 sky130_fd_sc_hd__clkbuf_2 output312 (.A(net312),
    .X(pcpi_rs1[15]));
 sky130_fd_sc_hd__clkbuf_2 output313 (.A(net313),
    .X(pcpi_rs1[16]));
 sky130_fd_sc_hd__clkbuf_2 output314 (.A(net314),
    .X(pcpi_rs1[17]));
 sky130_fd_sc_hd__clkbuf_2 output315 (.A(net315),
    .X(pcpi_rs1[18]));
 sky130_fd_sc_hd__clkbuf_2 output316 (.A(net316),
    .X(pcpi_rs1[19]));
 sky130_fd_sc_hd__clkbuf_2 output317 (.A(net317),
    .X(pcpi_rs1[1]));
 sky130_fd_sc_hd__clkbuf_2 output318 (.A(net318),
    .X(pcpi_rs1[20]));
 sky130_fd_sc_hd__clkbuf_2 output319 (.A(net319),
    .X(pcpi_rs1[21]));
 sky130_fd_sc_hd__clkbuf_2 output320 (.A(net320),
    .X(pcpi_rs1[22]));
 sky130_fd_sc_hd__clkbuf_2 output321 (.A(net321),
    .X(pcpi_rs1[23]));
 sky130_fd_sc_hd__clkbuf_2 output322 (.A(net322),
    .X(pcpi_rs1[24]));
 sky130_fd_sc_hd__clkbuf_2 output323 (.A(net323),
    .X(pcpi_rs1[25]));
 sky130_fd_sc_hd__clkbuf_2 output324 (.A(net324),
    .X(pcpi_rs1[26]));
 sky130_fd_sc_hd__clkbuf_2 output325 (.A(net325),
    .X(pcpi_rs1[27]));
 sky130_fd_sc_hd__clkbuf_2 output326 (.A(net326),
    .X(pcpi_rs1[28]));
 sky130_fd_sc_hd__clkbuf_2 output327 (.A(net327),
    .X(pcpi_rs1[29]));
 sky130_fd_sc_hd__clkbuf_2 output328 (.A(net328),
    .X(pcpi_rs1[2]));
 sky130_fd_sc_hd__clkbuf_2 output329 (.A(net329),
    .X(pcpi_rs1[30]));
 sky130_fd_sc_hd__clkbuf_2 output330 (.A(net330),
    .X(pcpi_rs1[31]));
 sky130_fd_sc_hd__clkbuf_2 output331 (.A(net331),
    .X(pcpi_rs1[3]));
 sky130_fd_sc_hd__clkbuf_2 output332 (.A(net332),
    .X(pcpi_rs1[4]));
 sky130_fd_sc_hd__clkbuf_2 output333 (.A(net333),
    .X(pcpi_rs1[5]));
 sky130_fd_sc_hd__clkbuf_2 output334 (.A(net334),
    .X(pcpi_rs1[6]));
 sky130_fd_sc_hd__clkbuf_2 output335 (.A(net335),
    .X(pcpi_rs1[7]));
 sky130_fd_sc_hd__clkbuf_2 output336 (.A(net336),
    .X(pcpi_rs1[8]));
 sky130_fd_sc_hd__clkbuf_2 output337 (.A(net337),
    .X(pcpi_rs1[9]));
 sky130_fd_sc_hd__clkbuf_2 output338 (.A(net338),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__clkbuf_2 output339 (.A(net339),
    .X(pcpi_rs2[10]));
 sky130_fd_sc_hd__clkbuf_2 output340 (.A(net340),
    .X(pcpi_rs2[11]));
 sky130_fd_sc_hd__clkbuf_2 output341 (.A(net341),
    .X(pcpi_rs2[12]));
 sky130_fd_sc_hd__clkbuf_2 output342 (.A(net342),
    .X(pcpi_rs2[13]));
 sky130_fd_sc_hd__clkbuf_2 output343 (.A(net343),
    .X(pcpi_rs2[14]));
 sky130_fd_sc_hd__clkbuf_2 output344 (.A(net344),
    .X(pcpi_rs2[15]));
 sky130_fd_sc_hd__clkbuf_2 output345 (.A(net345),
    .X(pcpi_rs2[16]));
 sky130_fd_sc_hd__clkbuf_2 output346 (.A(net346),
    .X(pcpi_rs2[17]));
 sky130_fd_sc_hd__clkbuf_2 output347 (.A(net347),
    .X(pcpi_rs2[18]));
 sky130_fd_sc_hd__clkbuf_2 output348 (.A(net348),
    .X(pcpi_rs2[19]));
 sky130_fd_sc_hd__clkbuf_2 output349 (.A(net349),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__clkbuf_2 output350 (.A(net350),
    .X(pcpi_rs2[20]));
 sky130_fd_sc_hd__clkbuf_2 output351 (.A(net351),
    .X(pcpi_rs2[21]));
 sky130_fd_sc_hd__clkbuf_2 output352 (.A(net352),
    .X(pcpi_rs2[22]));
 sky130_fd_sc_hd__clkbuf_2 output353 (.A(net353),
    .X(pcpi_rs2[23]));
 sky130_fd_sc_hd__clkbuf_2 output354 (.A(net354),
    .X(pcpi_rs2[24]));
 sky130_fd_sc_hd__clkbuf_2 output355 (.A(net355),
    .X(pcpi_rs2[25]));
 sky130_fd_sc_hd__clkbuf_2 output356 (.A(net356),
    .X(pcpi_rs2[26]));
 sky130_fd_sc_hd__clkbuf_2 output357 (.A(net357),
    .X(pcpi_rs2[27]));
 sky130_fd_sc_hd__clkbuf_2 output358 (.A(net358),
    .X(pcpi_rs2[28]));
 sky130_fd_sc_hd__clkbuf_2 output359 (.A(net359),
    .X(pcpi_rs2[29]));
 sky130_fd_sc_hd__clkbuf_2 output360 (.A(net360),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__clkbuf_2 output361 (.A(net361),
    .X(pcpi_rs2[30]));
 sky130_fd_sc_hd__clkbuf_2 output362 (.A(net362),
    .X(pcpi_rs2[31]));
 sky130_fd_sc_hd__clkbuf_2 output363 (.A(net363),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__clkbuf_2 output364 (.A(net364),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__clkbuf_2 output365 (.A(net365),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__clkbuf_2 output366 (.A(net366),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__clkbuf_2 output367 (.A(net367),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__clkbuf_2 output368 (.A(net368),
    .X(pcpi_rs2[8]));
 sky130_fd_sc_hd__clkbuf_2 output369 (.A(net369),
    .X(pcpi_rs2[9]));
 sky130_fd_sc_hd__clkbuf_2 output370 (.A(net370),
    .X(pcpi_valid));
 sky130_fd_sc_hd__clkbuf_2 output371 (.A(net371),
    .X(trace_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output372 (.A(net372),
    .X(trace_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output373 (.A(net373),
    .X(trace_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output374 (.A(net374),
    .X(trace_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output375 (.A(net375),
    .X(trace_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output376 (.A(net376),
    .X(trace_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output377 (.A(net377),
    .X(trace_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output378 (.A(net378),
    .X(trace_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output379 (.A(net379),
    .X(trace_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output380 (.A(net380),
    .X(trace_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output381 (.A(net381),
    .X(trace_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output382 (.A(net382),
    .X(trace_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output383 (.A(net383),
    .X(trace_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output384 (.A(net384),
    .X(trace_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output385 (.A(net385),
    .X(trace_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output386 (.A(net386),
    .X(trace_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output387 (.A(net387),
    .X(trace_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output388 (.A(net388),
    .X(trace_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output389 (.A(net389),
    .X(trace_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output390 (.A(net390),
    .X(trace_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output391 (.A(net391),
    .X(trace_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output392 (.A(net392),
    .X(trace_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output393 (.A(net393),
    .X(trace_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output394 (.A(net394),
    .X(trace_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output395 (.A(net395),
    .X(trace_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output396 (.A(net396),
    .X(trace_data[32]));
 sky130_fd_sc_hd__clkbuf_2 output397 (.A(net397),
    .X(trace_data[33]));
 sky130_fd_sc_hd__clkbuf_2 output398 (.A(net398),
    .X(trace_data[34]));
 sky130_fd_sc_hd__clkbuf_2 output399 (.A(net399),
    .X(trace_data[35]));
 sky130_fd_sc_hd__clkbuf_2 output400 (.A(net400),
    .X(trace_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output401 (.A(net401),
    .X(trace_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output402 (.A(net402),
    .X(trace_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output403 (.A(net403),
    .X(trace_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output404 (.A(net404),
    .X(trace_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output405 (.A(net405),
    .X(trace_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output406 (.A(net406),
    .X(trace_data[9]));
 sky130_fd_sc_hd__clkbuf_2 output407 (.A(net407),
    .X(trace_valid));
 sky130_fd_sc_hd__clkbuf_2 output408 (.A(net408),
    .X(trap));
 sky130_fd_sc_hd__buf_8 repeater409 (.A(_11309_),
    .X(net409));
 sky130_fd_sc_hd__buf_8 repeater410 (.A(_01208_),
    .X(net410));
 sky130_fd_sc_hd__buf_8 repeater411 (.A(_14356_),
    .X(net411));
 sky130_fd_sc_hd__buf_6 repeater412 (.A(_14355_),
    .X(net412));
 sky130_fd_sc_hd__buf_6 repeater413 (.A(_14939_),
    .X(net413));
 sky130_fd_sc_hd__buf_8 repeater414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__buf_8 repeater415 (.A(_00308_),
    .X(net415));
 sky130_fd_sc_hd__buf_8 repeater416 (.A(_20068_),
    .X(net416));
 sky130_fd_sc_hd__buf_8 repeater417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_8 repeater418 (.A(_20067_),
    .X(net418));
 sky130_fd_sc_hd__buf_8 repeater419 (.A(_20066_),
    .X(net419));
 sky130_fd_sc_hd__buf_8 repeater420 (.A(_20065_),
    .X(net420));
 sky130_fd_sc_hd__buf_4 repeater421 (.A(_19701_),
    .X(net421));
 sky130_fd_sc_hd__buf_6 repeater422 (.A(_19700_),
    .X(net422));
 sky130_fd_sc_hd__buf_4 repeater423 (.A(_19700_),
    .X(net423));
 sky130_fd_sc_hd__buf_6 repeater424 (.A(_19698_),
    .X(net424));
 sky130_fd_sc_hd__buf_8 repeater425 (.A(_18857_),
    .X(net425));
 sky130_fd_sc_hd__buf_8 repeater426 (.A(_19702_),
    .X(net426));
 sky130_fd_sc_hd__buf_6 repeater427 (.A(_18856_),
    .X(net427));
 sky130_fd_sc_hd__buf_12 repeater428 (.A(_02217_),
    .X(net428));
 sky130_fd_sc_hd__buf_8 repeater429 (.A(net431),
    .X(net429));
 sky130_fd_sc_hd__buf_8 repeater430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_8 repeater431 (.A(_02069_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_8 repeater432 (.A(_18832_),
    .X(net432));
 sky130_fd_sc_hd__buf_8 repeater433 (.A(_18810_),
    .X(net433));
 sky130_fd_sc_hd__buf_8 repeater434 (.A(_18805_),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_8 repeater435 (.A(net218),
    .X(net435));
 sky130_fd_sc_hd__buf_12 repeater436 (.A(_21107_),
    .X(net436));
 sky130_fd_sc_hd__buf_12 repeater437 (.A(mem_xfer),
    .X(net437));
 sky130_fd_sc_hd__buf_8 repeater438 (.A(_18816_),
    .X(net438));
 sky130_fd_sc_hd__buf_8 repeater439 (.A(_18788_),
    .X(net439));
 sky130_fd_sc_hd__buf_6 repeater440 (.A(_11336_),
    .X(net440));
 sky130_fd_sc_hd__buf_6 repeater441 (.A(_10404_),
    .X(net441));
 sky130_fd_sc_hd__buf_4 repeater442 (.A(_08243_),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_8 repeater443 (.A(_06529_),
    .X(net443));
 sky130_fd_sc_hd__buf_8 repeater444 (.A(_06369_),
    .X(net444));
 sky130_fd_sc_hd__buf_8 repeater445 (.A(_06297_),
    .X(net445));
 sky130_fd_sc_hd__buf_8 repeater446 (.A(_06248_),
    .X(net446));
 sky130_fd_sc_hd__buf_6 repeater447 (.A(_05978_),
    .X(net447));
 sky130_fd_sc_hd__buf_4 repeater448 (.A(_05633_),
    .X(net448));
 sky130_fd_sc_hd__buf_6 repeater449 (.A(_04840_),
    .X(net449));
 sky130_fd_sc_hd__buf_8 repeater450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_8 repeater451 (.A(_01683_),
    .X(net451));
 sky130_fd_sc_hd__buf_8 repeater452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_4 repeater453 (.A(_01683_),
    .X(net453));
 sky130_fd_sc_hd__buf_8 repeater454 (.A(_20150_),
    .X(net454));
 sky130_fd_sc_hd__buf_8 repeater455 (.A(_19900_),
    .X(net455));
 sky130_fd_sc_hd__buf_8 repeater456 (.A(_19891_),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_8 repeater457 (.A(_19878_),
    .X(net457));
 sky130_fd_sc_hd__buf_8 repeater458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_8 repeater459 (.A(_00309_),
    .X(net459));
 sky130_fd_sc_hd__buf_8 repeater460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_12 repeater461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_12 repeater462 (.A(_00368_),
    .X(net462));
 sky130_fd_sc_hd__buf_4 repeater463 (.A(_10987_),
    .X(net463));
 sky130_fd_sc_hd__buf_6 repeater464 (.A(_08614_),
    .X(net464));
 sky130_fd_sc_hd__buf_8 repeater465 (.A(_06446_),
    .X(net465));
 sky130_fd_sc_hd__buf_8 repeater466 (.A(_06310_),
    .X(net466));
 sky130_fd_sc_hd__buf_8 repeater467 (.A(_05512_),
    .X(net467));
 sky130_fd_sc_hd__buf_4 repeater468 (.A(_05502_),
    .X(net468));
 sky130_fd_sc_hd__buf_8 repeater469 (.A(_05217_),
    .X(net469));
 sky130_fd_sc_hd__buf_8 repeater470 (.A(_04837_),
    .X(net470));
 sky130_fd_sc_hd__buf_8 repeater471 (.A(_00292_),
    .X(net471));
 sky130_fd_sc_hd__buf_8 repeater472 (.A(_00292_),
    .X(net472));
 sky130_fd_sc_hd__buf_6 repeater473 (.A(_20129_),
    .X(net473));
 sky130_fd_sc_hd__buf_8 repeater474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_8 repeater475 (.A(net477),
    .X(net475));
 sky130_fd_sc_hd__buf_8 repeater476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_6 repeater477 (.A(_00301_),
    .X(net477));
 sky130_fd_sc_hd__buf_12 repeater478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__buf_12 repeater479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_8 repeater480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_12 repeater481 (.A(net488),
    .X(net481));
 sky130_fd_sc_hd__buf_8 repeater482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_12 repeater483 (.A(net485),
    .X(net483));
 sky130_fd_sc_hd__buf_8 repeater484 (.A(net485),
    .X(net484));
 sky130_fd_sc_hd__buf_12 repeater485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_12 repeater486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_12 repeater487 (.A(net489),
    .X(net487));
 sky130_fd_sc_hd__buf_8 repeater488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_8 repeater489 (.A(_00357_),
    .X(net489));
 sky130_fd_sc_hd__buf_12 repeater490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_12 repeater491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_12 repeater492 (.A(net497),
    .X(net492));
 sky130_fd_sc_hd__buf_8 repeater493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__buf_12 repeater494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__buf_12 repeater495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_12 repeater496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_12 repeater497 (.A(_00358_),
    .X(net497));
 sky130_fd_sc_hd__buf_12 repeater498 (.A(net500),
    .X(net498));
 sky130_fd_sc_hd__buf_12 repeater499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_12 repeater500 (.A(_00360_),
    .X(net500));
 sky130_fd_sc_hd__buf_12 repeater501 (.A(_00362_),
    .X(net501));
 sky130_fd_sc_hd__buf_12 repeater502 (.A(_00362_),
    .X(net502));
 sky130_fd_sc_hd__buf_8 repeater503 (.A(_12348_),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_8 repeater504 (.A(_11975_),
    .X(net504));
 sky130_fd_sc_hd__buf_6 repeater505 (.A(_06366_),
    .X(net505));
 sky130_fd_sc_hd__buf_6 repeater506 (.A(_01816_),
    .X(net506));
 sky130_fd_sc_hd__buf_8 repeater507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_8 repeater508 (.A(_01304_),
    .X(net508));
 sky130_fd_sc_hd__buf_8 repeater509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_8 repeater510 (.A(_00297_),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_16 repeater511 (.A(latched_store),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_16 repeater512 (.A(net226),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_16 repeater513 (.A(net225),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_16 repeater514 (.A(net222),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_16 repeater515 (.A(net211),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_16 repeater516 (.A(net200),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_16 repeater517 (.A(\cpu_state[3] ),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_16 repeater518 (.A(\cpu_state[2] ),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_16 repeater519 (.A(\pcpi_mul.shift_out ),
    .X(net519));
 sky130_fd_sc_hd__buf_8 repeater520 (.A(net7),
    .X(net520));
 sky130_fd_sc_hd__buf_8 repeater521 (.A(net65),
    .X(net521));
 sky130_fd_sc_hd__buf_8 repeater522 (.A(net60),
    .X(net522));
 sky130_fd_sc_hd__buf_8 repeater523 (.A(net56),
    .X(net523));
 sky130_fd_sc_hd__buf_8 repeater524 (.A(net45),
    .X(net524));
 sky130_fd_sc_hd__buf_8 repeater525 (.A(net44),
    .X(net525));
 sky130_fd_sc_hd__buf_8 repeater526 (.A(net43),
    .X(net526));
 sky130_fd_sc_hd__buf_8 repeater527 (.A(net39),
    .X(net527));
 sky130_fd_sc_hd__buf_8 repeater528 (.A(net36),
    .X(net528));
 sky130_fd_sc_hd__buf_8 repeater529 (.A(net30),
    .X(net529));
 sky130_fd_sc_hd__buf_8 repeater530 (.A(net21),
    .X(net530));
 sky130_fd_sc_hd__buf_8 repeater531 (.A(net20),
    .X(net531));
 sky130_fd_sc_hd__buf_8 repeater532 (.A(net2),
    .X(net532));
 sky130_fd_sc_hd__buf_8 repeater533 (.A(net13),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_opt_9_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_opt_8_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_opt_5_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_opt_6_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_opt_4_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_opt_0_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_0_1_clk (.A(clknet_2_0_0_clk),
    .X(clknet_2_0_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_1_1_clk (.A(clknet_2_1_0_clk),
    .X(clknet_2_1_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_2_1_clk (.A(clknet_2_2_0_clk),
    .X(clknet_2_2_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_3_1_clk (.A(clknet_2_3_0_clk),
    .X(clknet_2_3_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_0_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_1_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_2_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_3_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_4_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_5_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_6_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_7_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_0_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_3_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_4_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_5_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_6_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_7_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_8_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_9_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_10_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_11_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_12_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_13_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_14_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_15_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_16_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_17_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_18_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_19_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_20_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_21_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_22_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_23_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_24_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_25_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_26_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_27_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_28_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_29_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_30_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_31_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_clk (.A(clknet_5_1_0_clk),
    .X(clknet_opt_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_clk (.A(clknet_5_10_0_clk),
    .X(clknet_opt_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_clk (.A(clknet_5_10_0_clk),
    .X(clknet_opt_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_clk (.A(clknet_5_14_0_clk),
    .X(clknet_opt_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_clk (.A(clknet_5_15_0_clk),
    .X(clknet_opt_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_clk (.A(clknet_5_15_0_clk),
    .X(clknet_opt_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_clk (.A(clknet_5_21_0_clk),
    .X(clknet_opt_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_clk (.A(clknet_5_27_0_clk),
    .X(clknet_opt_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_9_clk (.A(clknet_5_31_0_clk),
    .X(clknet_opt_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_clk (.A(clknet_5_31_0_clk),
    .X(clknet_opt_10_clk));
endmodule
